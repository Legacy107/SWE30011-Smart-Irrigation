PK   ��VZ���=%  ;�    cirkitFile.json͝O��6�ſʆ�Z�@���6����ì��Cw�")�bʥ^��m����"�rW� %@��ef����L��D��վ�exh��~h~������-�w����ܾ���[}�>4�]�Ӿ��q��w����ۧ!Y_��9�5��ll�؂�$3y�ԅ)��l6�!���Yc�z�����H�4$f�F0�3H#�&3H#�&3H#�&3H#��3H#��3p����ϟv�á�z����d��u�U�N�kʒu��zkL1t�;Vws��u���Lb�|�jwZVV.J��ʮӮk���W�.�`�Z� ��R�<?�C8
@���h��hqG!����B���!�<S�C8
y��p�l-�(�S�Q�S�8���s�8����NqG��s����1�ܰdMպ��*1�b�dC�%��UI���������C+�Xy��p�-�(�9[�Q�s�8��%���l+�����s�8����lqG!����0+�����.-�о��֮mBά&Y�6��]�}ח�f]	sv*��c��}*��F���}�8������B�W�C8
y_!�(�}�8�i2y_!�(�}�8������B�W�C8
��|���s��z���o��4ͻ�J�+ʓ,���TQ�^o�23}���0C���9[�Q�s�8����lqG!������9[�Q�s�8����lqG!����B���!�ɣ|���s�8����NqG!ϝ��B�;�!LS�s�8����NqG!ϝ^�O���>ٷ����g�O��v�=��N~D�{~�#���d�����q��Vv(a�Lc��Y�vP:�鮾
�`�+{��JGX:�\��eX�t��s#�v9V;(a���]��JGX:ӔX�J�vP:�ҙ��jWa�����Ԡ�K�pT	�a�����X١t��]}I82"��"��������뇶Ch?6DvD�DX>����`����G`>~����`����{,����y�~`���#0����u�|��`��~�G`>^k�l\�|��U"�q������׷���,���Y��(Vh�-�a�i��w�T�Y�4^���z�|��P`����G`>^���z�|���g`����G`>^9��z�|��5`����G`>^���z�|��u��R���G`>^!
��z�|4�77�Z��J_����z|����D�4^���E6��I��'�,��x=2X?������WR���,��x8X?������W����,��x�=X?������+`�����G`>�u ��z�|��*`����G`>�/��?�|���`��kiЋi��#���?�|�� `����G`>�g��?�|��J,`����G3|sS�A�d�u��Xz�u����J��
��q���9��`���Ղ���]���|\����`�������]���|\[
���`���U��������]Ov=9��`��Ǖ����]���|\C���`������������|\��_�X>�q�=�~`���#0�
��X>��]���LH<�$�HHH2�j{Brͮ��_8'�a:'(@�^�霛 EzI�|���ِ}{�I���ߞJ��
��uYJ*E��[#�^��n�/�ӧ�m#O���+�&�A�LkqG���kN�B�ѻ��tXA_>-|{+Ho%�DҮe1�����Է�}���~���[�ۘ5�|��m�{���{�ƞ/�I�Va_/슼�2c�6_o������J3�%/oC�؁���{�0Fo��^`���#hdX�D�2YY�î�v��������l�:��Ռ����*����v"P ×C
d�f`�@�;(�a�!2l�0D�@������)JQ�"2l�0D�@f�u���ڸ���KܨHf4� &X�&X�FE2��1��7�8*�]:�	Ɍ����K�Hf�� ,ay���8*�gR@L�<nay���UWo�L�<��d�i ,�[XGE2�t�	��-,��"�q^���),��"�q����),��"q%����tk!,�#me�N���H\C���),��"q�,���<���5I`���<���8*�΀1��x��H\���g�<�G�v(!,��"��~,�g�<��ċ�aL�<���8*�\�1��x��H�����9,��"�JPl<���8*�X�1��x��H�����,��"�
0,��<�)~��ta <�<�{k�E��;hT�i��Q��j��
�i�	�Q��j�zK.ƨe.U`Z����	FVRau�KE�i�������A*�Nˢ`�`%V7FQ�uZ.��+���fZ@��+�����{|T��>+b���j�i�xT���^1�8�t�8.Zҡ�w�u�Ur]J�K�w���"�BK:������:�K��th��ymu�
-����:��0Zҡ�5:��81Zҡ�:��1Zҡ�5%:��82Zҡ�1:��2Zҡ�5>:t|�
-�К��Hmu|�
�_4�0����V鉘O��S��c:���2Zҡ�5p:���2Zҡ�|:���2Zҡ�5�:���2Zҡ嵕:���2Zҡ�5�:���2Zҡ嵮:���2Zҡ�5�:/&��2Zҡ5'Š����2Z�"6�}:_����Z�/S���:�*�������/Ku|Y���ThI�����h���ThI��k�h���ThI��k%�h���ThI��k>�h���ThI��kW�h���ThI��kp�h���2Zҡ�Z":���2Zҡ�(:���2Zҡ��.:���2Zҡ�5:�*�$SZJ���2_���2Zҡ�A:���2Zҡ��G:���2Zҡ5'{�"���e*��F����馨(mu|�-bn\��kj�h���2Zҡ��`:���2Zҡ�g:���2Zҡ�Zm:���2Zҡ�s:���2Zҡ��y:�*U�P*���r_���2Zҡ�Z�:���2Zҡ嚌:���2Zҡ�ڒ:���2Zҡ��*�:�L��th�֧��:�L��th�f���:�L���h_���z����d��u�U�N�kʒu��zkL1t�qf")2
���EF9V��v�}�Rn�4��*)�.O��s�"jS���ۼ����2KP��KP�����=^��m��vmr$Y�6�'�Sh��]_��u5��+Od����EF��t	��^�FA��/Ti���PW92�B%��(5�#�d��QP��:�Q
ȕ^�����_��,�+�mu�Ƌi����%��0�Lfaۃ�0����nlL^��66�/m$��/v�aa0YxiS��0�V���hlL+>n��obӊ��ьs�����*1�b�dC��بJ�v0n�W�`���s�E�8~�b_��_�0�a�<�ðz��K��M(�W>O�}{��/~
P 3*!2��"P 3�O!D�@f�B�@��8n���q!2�xB
dFo !2�π���g��H\�ƥmX�&X�FE2Gk�a��n�%oT$s4�&X�&XGE2G;�a��p�%qT$s4�&X��<��d�S &��7 ��q��H�8Ӂa��q��H�8�a��q��H�8;�a��q��H�8o���<���8*W+�1�fRpS)�<���8*W��1��x
��H\����),��"q�,�g�<���U`L�<���8*W�1���q��<���8*�ކ1��x��H�Z���,��"��TأX�ay�WC`y<��qT$^}c�=��=ބ����Q�x��	��sXGE�U90&X/`y�W���`y����H�+:�C�ǅ����J*���V��u�`%V�x+��Q��j��
�i���@]5XI���.]��4XI�Ս�Tt��6@�`%V7FQ��+� Q@��TXM�Uk@G��J*���*5��u�`%V�xU�Q��j��
+��ct�
-����:�*�.%ۥ�H�x���R�%Z~�\G[��BK:��μ��:L��th��mu\�
-���mu��
-���Zmuܘ
-���mu�
-����mu\�
-����:�L��thy����:�L��thy͕��JOĔ���2��ˬ�/S�%Z^����/S�%Z^˧���/S�%Z^�����/S�%Z^[����/S�%Z^#����/S�%Z^몣��/S�%Z^���b��/S�%Z^{����/S�%Z^C����/S�%Z^����ۊJ�+���TǗ�:�L��thym���:�L��th�ƀ��:�L��th�V���:�L��th�惎�:�L��th�v���:�L��th������/S�%Z�%����/S�%Z������/S�%Z����/S�%Z�Q����J2��d:�,��e��/S�%Z�����/S�%Z�}����/S�%Z�ᤣ��/S�%Z�E����/S�%Z����m���ThI��k��h���ThI��k��h���ThI��k��h���ThI��k��h���ThI��k��h�T�C�̇�/�u|Y���ThI��k�h���ThI��k2�h���ThI��kK�h���ThI��kd�h[��2Zҡ�Z�:���2Zҡ嚥:���2Z
�}�*�ꁪ���M��IV�:Y�)K����1���K�0GFY�Me���K�r��y�VIQwy��@�P���L�����ґQ.���(Q��ik�6!'@��k��y;��i��e�YW��_��/
���E��#wn��KP�����i���e�j|d��:�Q*�GFY��e��yd��z屭�x1�wi���0����-plL^�|76�/mqӊ�6�����V���jlL+^��46�/�ӊ����u1�xi�˗0n�����J̦�$ِv<6����F�U7�ˣ��(��7ԗ;����nw��7����[J�V�����t�vC�l�ݾ�����	�/"�4�3�pw=I!#�X��@k�$~��R��F&CtA}���� i�m�.˓b�L]f�:���$mZ֖Ҷ6T���肸n\��$�v�m�~��E��¦9-����iE(��~7D��"wK���8u}K�"����7p>I�����s��$j��|�[�L��)]�4?��k����[#3¯�%_OV��$��T����<�-�=��D���x�8���oZ�]´�4IR��IH{�s����#�i^L�m�bvӯ�t��7�2a3�b�>-)�tG���Zd��2�J���T��Ҿ�\#����8 �*I��������8��!p��[t�g'p}H���Ç?����ϻ_��i����w��<���f�_��?���O�@��g��ճ9��!�?���@?\J+7y\!'B?�8Kt��Ӧsk���&OUn����g�(�^��S9����,�Mɉ�O��D�C3����A��B!~Z���>4�P���ǘr��O�"�i��}���4L��>T\����qc|�[w��vj/�c�����B�G��~0�H��._�۸wD�Y���4��f�>�����O�Mg�~t�����ݦ�����x�6���BlPZH_R3�(-�o��%��!�T��;7�^�o��a���hn���'�~'��'�n'�C��	}K;�s�k���}09��09��0=c>gj��WՖ��M^�A��~���>q�oo�B���.�2�u����������ۯ���l�ћîy�����_�j�z�,[�C����B���f��$��0c�(!�8��L	)�!�X�JH!a�*WB
aN�=l1c�,!�8��n	)�!̱h�4�!�)"��)�<�9��r R*r�<�9V>�r �*�<�9�^�r�c�c�6) � ��c���<�9֟�r ����) �Z@>c��DH4id���X��j�U�k�I9 ��ҫ<�9V�r ҫ�Wys�k(5����ҫ<���r��GL ����B,@zcL�J! ��c8@���p�l+��8 �V�q ��<�i2@���p�l+��{�8 �6d[y����f�|:Ƙ�� ��c�� @z� �U��3p �kH���M.��^s@z����W���ҫ<o�	� Ws@>����"�|��<oC� ���O�1x{;  ��|�ǈߒ����g�(�We�s��7�����v9�Ńȉ��^S�^o'C\<�~X>�:�y�^G3����PNo7y�����Ϲ�~ގ��ߋ�#0�}���v��^,���(������b��go�w\<�~X>�i�Dd<�~ߤ�. ���ۻ"'�ϫu�]QV~?=�F�0!�	��N��p��,h�Bh�Bh�&$4!�S���U���&������
��Є�.3ZC�g����Fk��-`BB�;�h��LHhBsR�	�!ڿ�	��V��,�6-`BB���6ڧ�		Mh�2vЀ�>�'�<�n��\R���p� �"���]�E�0!�	y�ZC������5D�0!�	y�ZC�����j�5D�0!�	�W�!�ŀ	�I�T��h&�k����@���b���&4'%1�]��/��=��
�]L�v1>�D��Jᯍ����8�v1��1�]����5D�0!�	y1ZC�����@�5D�0!�	y�6ZC�������5D�0!�	y�<X��b���&�%�h�.LHhB.W��m[���&�Rh�>LHhB.�������S2�O��>LHhB�ǁ��S���&4��Ѐ�>LhN��h��)`Bo~R�m���D�K��->��=�BBsu��9�ŀ		Mȕu��]��Є\�!�ŀ		M����]��Є\�	�!�ŀ		Mȕ���W�×�]L�v19�ŀ		M����]��Є\}�!�ŀ		Mȕ���m��Є\��a��)`BBr�:��h�&$4!W�Ck��)`B�D���$�U}_'�<����u�^S���u�[c����-��V�G~��-���Y?����������R��|R�~��kaGo�|~��}����;���%�7�?��i�~�^=���:������ G�?���d�g�q�����'F�� G�_g��p^���&n���J3w�Br�7s;/䮰x^=�� ���>@�h���bH۩��^l qZ�b��I󬿋\l i���m� m��O�$�l��b;Oi;��{	��}몯��l�M�iǣ�*)����a_u���-)nf���}�����՗��K�m�[λ����|�H��݊"s�Շ�UȈ�;)d�xz��*�C.��݊���ѱ���ǜ<�/�(�_Ƃ�7 >��p��O >��v��gX>���ϰ|��3,�a����pM��\��X�z=/��p�Ը\(o��N�~)2��	Ξ�]�ɹęJƏ�oI�4�"��KBg8a)��̥�[A�0�:�Xj�ה�_�0:��7x���wh&qV2Udg�M�p�P�n��j[����Y!���B�[�]h���)����5��u�pL���v�O�ԗ��dt��v�3A2�Kp�\��2�uM��.�Á���W)_� ï��]�<��(�^�?�ÿ�8�O��G��(}�(�?ʞ?�����r������������������~���#������\������i�g=���x���#�!��w�����U��>lv������*�����{���.�}s�Ui���!/��as����������u�������O���Fk���?�%�P�����''�C�3�7z������������7�����+�o�w���7y�v��?���a����v}?|��~�ߧ�~p>��~��?�O��;<��9�ׇ�������� �cq�����9)��y�V6�CP{GY�&ͩ6i}�'u�2��\�UV�͊!I���U�'i;���L[m��0ۇ�C���	��w��~�^{[�?}<��v�}w?<_�w��o�;����]A�˿��MV��S��0�������S���c�?��zc�2�DN婳7U���z�[�UY���[6Ϟ��:뢫�/���Y�Qf���$��զ���|�T� /?U��}~��!�9�we�;uj;��r�x�j���䕵�-MQ�-��*�ܟ���,-���u+�����~�un����j^7�)�օ����4�֪/7��⦔�kcUV�im�mPUT�ĵ2��Җ�.;���ʉ��-]�r:UoJk���}�ur�Z�m�t�np:m։�L��4��tݥk;�)h�l���'O�t�����x�wwI��7��'E��Iuz�u�-*��e�2�?A�˾�>��I<��k4�]>����mǦ�:�L��{�$�:vIk�:����˼�2��M�����c�6�md��d]��(�Y�������IZ.}b�1K�P�t^��A6aN�~2�^>��9_��3+MU�����Nؤ�O�E��YZ,fϜg�ɗ�gk�h�p\Y�W�ˊ�UZ80��)0�LY8����^�Z8�og��n�@�.�5���6:sإl��a��ЏY��sIq�@�1��+�h��-������Cج~Cy=������s��n�2�J��:=���/�Zm�q�����������>��K��lc~ﺤ�������տ~���~u���������o�����Q�`�C?J�Xe�o?��Du��C���n�p��=|c�������7?�?�}�#���;�߱Ox���W�����;,ͧ�}��~�ŵ����qcڳ���'Sg�x샪KW��.y|Z'�����9��B�����^]�,�g/�䰒�[��>�07���7��'����Bn�
U�X�:����չÊ���|c��HC;��ʎ$ؑ��F7:�!���n���Ĕ9�r�r�>�_nB_�����j�Ǟ�ܧ�-�&��9=,M�	j���ԛn�X�׳��8$M�}]5�yзL��EP;=,�k�es	{5F��[#Xe�ea�:9��?*����FP��-:t#8gV�_GRl:g�W5�2d<:9�ԩ�$������q�����j[�fh*K���2��7��;ji��� nY��Vq�����a�edi�(crTB��&���*���e�	{�S��g�VYsY��}����l:�[��܉w����q���p��o+����F6�i'����ǖ�G��ڨ)������^9��l3��FQ�� �]qT�DYg��ހ;f^�^7��Tl�y�`�l�o�-u��Bm�-/o�� ��d^��dr�������^|�|\� 3��[��$쵝D+���Íl>����;� ��$a^���ab+�bˇ�e�ey��/�b���^�+�u*�Z��Y�*�ѿ�a+���{�@+�zG���n�/�/7wT6?%U]q��Q[.�m:��c�Vdә��m:T�4
y��W�4��WJ����o������皌�5=�������{�����u����Ϗ��>|Y}�PK   ��V5���� � /   images/1198b7a7-cbce-4bfb-9393-e70c622bc3b2.pngt{T�����������	�,�݂��E��`	��%$����o��{��|�;g����骮����T��I�  ���� �  �eQ�aW⏻�  LG[))5))j5W'k[+ @>:]EOs�8� %)	
�*�ցF����ؕ�MOB��&�͘�Ȱ-�\FW�p=�)��-��	[9�~��r8��/�N�N��G��cA#y�(�q�h:���&���8�q��I�p����Kpɣ�
zuuꀑ���#���
=����,B�!q(�l����� Uv@p9�@�9��<��#(J���+��ƪ�#y�B����K /K�82h�r��g!In���üS3�7jԣ�$�����9#��`�'��u
O���Y�o\���t�(�Zy���{q��.zqU��>d�J5R��CT�':G%�H��K�q	�3��84��G a����m"鹥��8������u�z�S��"�Hȋ#b����T�:��X��$��q���t�F>�늋���p]�&8�-
lD�d�������hf\M�,��rR�pul��4�xZ�(�G6�N$�9q#��o�z�l��#�t&|��_e�֥�Nz��̛���)��31<�R[�c��ZZ#��a�J��XL"�� M�(H�����$o~�<p��0Δt��k���B����9�h��nN��.#��g%r㊋4O��+�<A�m�n�e���1ɐi����!bF�1�VȬ�D!��9��: �§�$���X]{4��%�º�����Sz����I�)��q��=t���u��|�>�"�Da�~�oj.�:�H����I��9Ĺy]iɏ+��*�,ܳ���Ce�JzJdG=�"I\K;v��>d��#�zv��rn0>��������`�P�L�m���؄��G�"\���%�0аb��������R} [P��
:�����]�s�,�o[+5�� ѓҾ�`߻W�s�	�s����j� iI���	
S�QW�R���1j�ebj��ZǨP� �����I�����-������nT�p�K��-qaе��;�D3(�yʩ5���ݳ��3���U��p��]�#��!ꉉ$A>P��-�bl���U�MM�<��&��l���#���=|i�3��ұJ]���(��:�*Ԍ�����-��FE+|�ޏ�Z�O��Ȍ�I�}?m�<rJ|� 7BVbk��N	�`0��
�v��&���2u��Ǣ�r4���,&�xi��S0��KvI��k#����"Fh�G#B@��9@s�������b_=3k�H�jd���[��*����K=k��}�'�7��$Ʊ���qN)XCd���Q�{�$���3�d�%��&5�(��g�w��U���[F��ˏ��}�?�o�m)�Jw�l.o�W�٘�9#�*�G���ˣ馍���IP5�ɪ�X�ix��X=�B��T«���ѡ�a�M�MW*�s��b:W&7�4����K��;�K��ǽ��ʠ�=5�r;!m�7�ޕ.�v~��5��Ik�����+���!sγ��^k{-�����G���YK[(�w�i����j��o��v��+�BE�U�9�D��
��E_9������z%䟇$�讲'Rj�(�3Q<Y�TVP굇���C�U��c��Ǣ�߅���e�e����>t��݅�������
�8f��>�t~݌�����5d�f^;����(ae�i�O��^�99L=w��XY�,�5r��b�̘�a�Dx��.̥��}��@�@C)�~��r��2����n%�!wq�mN��NoV���k�8Y�����y�%C����퓽�4�����b�?*�Z}ز%�d�z��S]Ys��Z�5+��e֦feq�g�<[cE�����h{}�����][��|�d��p��ǉ3������4�(�LŢ��w"nb9��t�^�+�{���N�1���d�����d[Z�8ᳪ�H��Qό�bwY��l�J�2]�|�������M�MsG	G���GM";�"ľ����gi��ޞ>o}��ߝ��XpgpM��������]�^0�}Nu�t츲]�NC։�q~�7q���羂����o]��"�dj/O���ITʹ'/G���~��m��a	�_���;b���*�.J�K�H�F��~AǮ�>D;G͡�%WAM�4�L��]s��3��U�Ѡ%����q�J�卓��{��۸ѣQ�����\��R��<r?`�2]�k`��C�M�Ex4Z�2=2=�b{�e���¬���7�����-��x��x�}�-K��2�Yr�����ЦU���.���FY��xXr9܂��ѕ�r�ڲ��`�f,~M�ՏG0�����aYY1�:��Kq�Q����V��}��&W�f��J��汳�����>d�m<M��N&����Oxu	��v)�%�?�R�-����i?
[F9�Ww�Hg�F7Ň���Ht3SD��Z��5����W�L�;�7��^���=�-����f�������\>�9Ñ����q��&�e�s���l\o�lz6
z+9f�>��9���'��͛����e2y0��>��7m�Nr<���~�j�?����A��UGc��S�O�X1c^k�C����A5YͿ���~I�r��bK}�r�z���ڧ���2@�϶|H����cǗ�����6<ZScf`���e�+^��_�����If��!�O�֍Q�Ӊ��6mm�C��jҚ�^�
+n>N'�w�e�5���G(�[�&�C���=�Ƥx���[׸��5�k����ͩ�ҭ�+�9��O�y�e��O=غ	�xT�Q�O�}D��H٤����z0l_���%/A$�Hi'+��M��m��ȱ��������$���8ϿO��&��T4����3qS�
|xӝN��9�e�������L���RׂKl���a���c���6�m�5�ယ{+�8*�'���N���0��bo�ݯ_��2�3��|e�����k�?��4�9б���0g�yEEf��qw9�-n�7p�����(�a�fm1/����w���U����kz*L񃻡�+͑2� M�T������'�g�OO�h�#7�ݫ��z�w@��>ߤ>���'����Fc��w�A������8X�^�����C���p##eI�jiai)�U}%�s�������v||\up�\����7h]W����w�i �i��&4�v�颍<�A�hu�0��}�i�? 1Vz
��� X�G
@���`��ʲpL ��ex  �����*�~I�:�爐@���a�7�߭����e�t�ДRP�5-\����N��W9��h��o�  b�?;���	�׬����������;3K's+�w��/�-+��r7��~���&�-J����2'��&���4z�j�RN�V�|\\4b����"���BҲ��;���;qrzyyqx�p8��p�������f��`w�qt7�fwt���&�������������#��s3s'wQ�����σ��m��I�n�l��j8_spq���n�窐�����[i�w0���!�+�-����������zn���S���v�r�rz�v�u������� 8��$�3��,�.������:h@`j$��VՂ���Up��?L�a;����  (HKhy����>u-��#�'���2Ӕ��Ҙ�M5d��v��c!	�y�o���D��{��������a�q��ω���zy������;k3c�?��V%Ť���ʾ���KWSA)��EH�T�(���=�h��J��[n
��r�0���1�_���|�t[�#ɾI��T��+�E���kN1]��r\agtЛ*�,c;��mUk.�"a��Z�Ve��'��o����k�R�y����T/�Y���z%���Q�1�*�D;HKE�)�vB��PL���kه�,`o+�L�q���~�Nk����D�?�Z%p�(� \���% Q�8Ւ��r{#��:|y��� {�!�X�kT��S�P�3�� �oҐ���ğ̞q�T��@��2��SE��N/]�07v�^���v��^5�C��4Hw~ ȑNs�ޒ�=I�v��y�#AQ8<6^�t�C�GF:��D����;ʜP��9n ��$���A˺y���D��eWȾ�'��FNA�����9�!�L1�X��X�\�iA/
2���?�o���5u./�8���C�d�s�C_zZ՞$L�W�&�a�
��c���C \d��,g�C	*#*�?i�"�d2��dM%$"C"X�����7�.�{�ie���a����p��5�%�x��3�:d k9�G����UT+�<;�2��[�KXE��F�(iS"��K�j�'T�f[�5<�+��A�Z�ԢdC�T'�u��@_�0���k�}�{zsd"�WDޖx2)������P�7��^vv ���{�.Y��\��U	��;m�W�����BFn�����m���%�@�е\.p�,a"�zߛ��cJy�8�F����K-� Ҙ�*%�]�Y �(�L8Ƙi@/�� �N��4�q�9�PZ�_�R���xE��fv���c��*}����,�e��_vBs�Q�<�����>a���K���ٞ�
!�Eb8g�ԡY��,�]T###ᒽhֵ�k�@�@4�����
�Iښ��J����a����a��vkf���YM6�:��`tbm49��co=Pf�����4TP�)�4��RN_.�ڂ�c��t����:E-9SNi����(��8�*�X�O}�G��	�`ok���p��]n]��%ٕx,��J�c�*E�&H.EA���=ȃ,���ɀ��aS;��i$P�$5J��5h���Kb'�����EX���c�R�n�v���(��> 		��64��)U��M��V�Rz,��,8�H�=����F\�>�v�
EE�O����1CՄҜH~sŗ�F���e|�Á��a�#+�U���������6V$F�΄G����DD���^;��3��4g���y�Eæ}�}AW_���c��:zl��VMx�Oڪ<�.�}���gV��|d:������!��@v .NVU��N�CGV5{,8�[��� �ZM��X�\���ػQk��K촳�GiF�t{�w#�Fx^�A�d�w��e_����_�|ݱ������1qa�����KR��U��#���ӟ�1�Y�G�L���bl����=����UvU"O���خ6-��`��[k�rr:� �����ܗ�;�eٻ]?�y��*��b�M݃���.�Wq�a�����Խ���)�<�q5m���V���_�k1��q�huF�����0{zb�������A��O9�����7!1#����3�a�ubE����w�EBd�5M�J�������������ImX>z%/Gk|���kv�h:���{����R����I�Y���y�>�̼��N�
q�����Yn��x!#��=ܘK�1pZD� ����-'���1:��(g���m�\P�L;w=�� )���7U]^t>�C�u'��:�lb�>S��>��)�M��"�Վi�u;�4p4p6^T_�~��m���*a�Q\\���~�:d"O��R��Q��td���s�s�,�M�z�|C`��������8y�ߒ0� W� �'����%ľ  e��t$F�y�.�/���E�D��l�xE�O��
�tC8��?!�
g�S���;�B��|Yа#�	�<�@�V�Ba=�sj.�Pw� �JA.�rͩ�Y�G(�@����GVV�H�_���u����Z�]&A�^ڶ&�G���C�fO���8�̋�O���II���2�+�>�>_��?^-�׾�"�ܦ��.���Y���{C���
����� ��+�\��NA����*���;�ֺ}���+���@�1�R3�)$��\���ޛߒ2�Ӵ���.n��.���chC�%�jс�01i�F��0��\�h��_'�np�jX��Σ;��{iQ��B�۹:�S�Q�NTO����b��T�.L�I?\O�R�Í���ܸ�>l|�s�go��n߆J�p�{�4�Df��]u�;uH�|r`u~Ba �������p��b����I+|��$�����"yD����H�'��w�:��|1Y<��7�����f��>'=������[����ƚ��cV~x!s�R�:`�֌��D�`[�󠢬 ������U(���x��}�1�d,��\�����|�m�I�:����)o+'ym���֖���L�d=��7�����VD`M'x`�n
ل7�UK����q�)��,ҳ)D&���T\}�gYK�}�>B�rC��"	�KH��F�"J��>�o�L��nU�C���5O�m`�ƻ�lGJ�BU̸7�r�V�2yb������0�J�(GfA:K�6�#�������N����'��O4�[,��vߟ��Ѻ�&��a�Fn��f8�^"�8Q�p�0���W%��������5�XG1�-�:��	�S˕>x���)�ӬUNU[�	0N�Ib�آ�)v�����~SDܘ�#��9������52~��|������)�6��΀6b�YMyo\�s�����@b�J.�*�E��0���78e�8���ϻ��ŷ�֯��z��<�Y�w����;�LvK=�Ҥj�Q�iGD�\���a����r! ��E�[�,�3[#l�K��'���I��w���� (��wM�Gx��::Ȫ��qSV�k����n<%%%z1�Ɏ[�z��Y���!�r �	������V���]q����,"	�6ϐ�[5]P�����j�q.GG����SIii�/��WmX���I�L!wI�ں]�&�𡄊�Ʊ����`�n�� .�Ɵ�Wls!*��!TX��)�� U��'N�ͧ�97Ԛ�H$�?d%�iI��hnW^�bw>��~��N3CC�����Y؝�s2������t�@a�]Xd�M���r񭤎��9E��`y�B�4͉�A"��c猴�_�,܍0�@�(t�Uw�]���AT`\
�k�BOfV��>ժ͊�ڠ�B�B-���y�w �ףl����͎���re��|V����l�Y�~V�{�k�n����Cm�I�Y�7��~�rJ7;�a�031�dΆ���|]y�w}I�7�J���W$�С�����ã�#��f��!����ݎ������$���s��>�-�󨎼�G��g�j:^��>0(���wY�������rӭǞ��P±z7@����
�VY��T�����էڭ�G�o[]_>�x�����f��O��~�km+��c��W����ϯ��k�S8ތ4<tg����W���%q{ �kJE��
G�FP�������R����(���5J���<-��|4��=�E�H�״�BVB�t�j�Ԫ$4��K�5$�������H���H�1L����f�;�^�/<��+\�~��g	�8򵤠�
���
�� ��iw�d(��ޅ�8QA����ʠ�_M\^��f[�`W������������jKŤ�6�*uY�i�������9n�i�-�c9�P"!��OA��Q��>�2U���O�Y��+�������Or:��[a�Ndʪe�����ż�t��J^D�C�r�(>YPW$��E��koҠ��=���I[��=�`<$PVp<�xs�� Q�َ��u��_�d�Ԥ$ O�dpl��*<i�%���@��KLy�G,�ɳ.n�H0�ǿ@��,�MIU��9/F$�D~9���D�'�E��:lrM>�ox�f�P��$?���M*��1��t��H��-��~H�7�P�t�Y9��j;=ۗ�\��Qx���an�a$��'j�Lo lpD��򦄹9���a1 "O3�@��
1�ͷ��Í���������J��v^�n��u��v~@»=,^Qd7����+���\wk����0��R:�_��iKY�ey����6��,����ǻ__�������~~�3	P>/���=�l=��O�E=��}L���.�s�{%Zʵ����9��MQB�%}�0�-�|�o�Y�ll�>fÏg�6�٬��=���zS��A�̐��#eoI�.F��_A���22lo�1���ޠ�0C7�1	��}��?��Loh��91R/�Aؾ(��W���L1�7g[�k6�0������&��]�\�έ�.�8�C��T^،��z�q��|9�R����@ݜ��R}�k_��=��x�P�L�wŏ�^o��o,2>`��{]kev|}u$�bF7���ӎzq|��Z$6E(
e;���&;��g�,O�S�(g$�$kfQS��]��B9E��M� o���1\�NM�{���*9�>�ι#�n1�K�I'�:�`d3��hȵSy�TA����71D������yyy�1�6��#������e�Y��r^�}z��|7W����kǠ���ʠʬY�T�+�4�
���؋oL��a��������|���L�;��Z�ϵ�,�];&��D.��UAA�M�?�"h�=#'gT�6[JR��p����������[:0::z$�%e���i����D^Q�:E.�s8��6"$��qZ�V=����SF^J
:��Ӏlɕ]�<V&Z�I/FavH��`�Y�\�3�Q�M��|�6�^#8���gFzz$�/�}��|�DVVV��O��ϕ��p`4��@�6ʑ��2�<x,�9��÷��[��躢w�6�ܟ�5{��c��� �I��L`C��FXG�0M��w��T��º5u'���N�������!vd���W����	��	�:�'��N����Q�?�b��r�PS����:�]�߰a�o$���^* ܺ?
�+�ɟ��~sC){���g����Ք��44qQ��e���h�k�k�����wx"�O�(���Vc��xe@%o``D�R'd �@)�ٗ��r�Lo�U�������*����j�T���j�������E�F𞫪+�cb��>�����9W�[���l+s���\�@����*H{�!���;���q������f�,`�GU�Y�?<؞@�nn�O%v�ʋ3S���J��z�%�a��Lş|����G�����\Y�%Gk�L��0ccٹ���Q2����W�|��,׫7�'k|�fb�V�G6D��E�7|?ݑ��� �:�?�ì2�z1j^�'�Yȹ��6�
.�bcb\���ӪXd��[���s�K�Cu�J���
�s\By�^���nxxx^��N�"L���׭�j4��1��=�R����S�t�N�,�=?!�պ���C�%�5 \`�Z�G{�Z你h�~^���E1w$NU쩋���m:{"��6�JGO�������y/�啕��W�	:7CH�j"M��4���N�H��4oN�z�]5��E���!��y�o�V�PZ�⧎��Y�`�M�/x;����E)@��>�����]�u��;�RR�������f��0!��ܼ��^.��(B�TX\2%���ȗ��*sc�h(YYxȀ꽱7����"XH�m��3�@�fj6��/&]���S��`8�o�kw7�!���/p&��T���PS��_��y�$��X�\r�qlU����/ X��,��k����?��,pd�����(�p��\K'�u���kޠA*�ӳF/�H~��>�Mu�<�&;�p�SH\>svD<��4I�D=�6w���A��^�e���q�Y����<��Ҩ�V,���ɵD���$˟d=��>j����Y�*/������fd�`Ѻ��ʫzT��i����F��������{c�w�<ȝ�%����<o@�_���v!���0�M���������^a���UԀ���*��]J"VC�6ږ�!�Z��ѡ'�j�Zb�yϭ�&~�����1�a>*��z���e���N���c��5M��M�<s�vy����8q�CT����KmS*�!~��
��v�	\R?ۗ�$�#S��"i��	X�B�v���ɗ�?��V��Z�⃫mU<�ڢɶ�]S�P��W�AlHU���m�\�I ")"YG*�x.�:�8U$U�!��j�(�הF�<<߭���)�X8x�)dp���t�r�q�Fqg�nv�o�� �ޟ�ҚĖ��Xe�j��m{ħ���U�����
'��7��$TT��0�ٙ�ק�;��TN�Q�lz��tj�^:t�hLo�Ҡ�Ӄ���,��Bf�QE�v�
7��ZO�����4����)w�@�MI������J3�d�J\(�
4n�[��Dg*~/-�g����.ȩц�ìm:��&�n,� �܇�cD�|��~&�Z��V"r����;��[�95y>	�'�i-n�V��a��y�k�O#��ԭz����;������?�b��7�6�0���ʠ�}r-N��?�\���D���RFֺ������h�c�lt���4���j}GЧ����v��N�2 3B8���P\��*�)��JC-�+���Pz��N�fcv
j����~��@M|�y���ǂnQ�yQ*0�h;�
����~�G�_$K���05dӢ��'nzP��E u4/��H<k�� ��	i���l�b��/,l@��D_����$���ø���س�[:�~�v����?t�v1��{�n�Q�
�	
�?|>h�4�9�>��$�.V���= ����ס�Z9xL/*f�!�Z�x��@jҼ�f٭4P����ᄜJ��]��������\��F]�B:Ȩ�A�fWx	)� ��܈���um�Gy��j�
�pp8��Ħ��8$"ܓ��}�Zka�4��ZͦTb��)N�4W�ki�z���,Z�W���0��X����%��.w.}�V(&||��D$S'%L7���}�A�G��R�i}ZKN��ŀ����H���V�+'��rr(^�X=\h��[ߚ���Rؑ�fi�/l�̈́,7�m���eb��.l���m���I���Z��Q�)���y$����8ʭ�}.Nw�K����M%��"%��#`H��e~	Fv�F�}�$E�����߫��򸦷W�3�r��<B�:��_�U��ߢV�%��cl��ն�~JPO(�Z�ӂ=�J7�I��Ic�Y�.��`2��L���`���4������u"H�R���}ٰo�`^��]���T�(Џ�j$+�eW�d?j-��xm��S��g��17�b?Ӣ��F-�gF�^jM��΄U�TD�H�D��׫��Q�yѰ�m�׆�f!���	�%����U�v��S���V+�d=�^:(b���e~CC6��<�N]\p�� XgKI��0ȅI��^\T$Z���&e�6K.3=���[>J�$F_�ykkK�Y]�=	�IM{��K�*1�3.�
�����-�%e(�j�t\����^�����x�)����A���z�R��.���j8��`��s�
E�G��L���9~����q����٧�l �(@�Ġ7~N�E ��W$���]g��ژ`gtZʰ�Zy�ўħ��LI��wR���m�c򏷫a8�ؼ�<͔i�0��E�׻���_h��� ����[L롶�bD��� �L���^��W�P�����['�52bWniJ�$w�@j��ƆJ(� N°jiۛ�E�Smnw�����(��Q�ld�q���)a�n?��1�N����3u���l oYSA�C���/�fb`J������sj)�r~B�Е�N��~r��LRA�a6���-a ���<; ӎ�׋�.MTīL}����ǌ��F�ڿ��ս����>�P�u#�1)T���O�,%e�:��ՠ�ISK4]h�rc���\=�646t�Q���ג!k�j�K�¥Z|�]�����c�R�U��J����8�������$`�/7�^4ZsO�{�c���rZ|Y8W�M��Դ�M����Γ|&����D�ϧ=ȟ��(77�=���)l.��黦�6g����%�"��G�E�Ǜ�.ȗv�=Y&!�����J�6v�3�d3(#��vzt�)jGa��eTU�8���ꚑS�fGTꘇdq��*���"����~�G x!E~�ͅ���H����%��[@��@9�ZU�5��YfW�z$�a���D@1{����>f?}^�Y1�!�L2�n�XC?Qÿ��P�[��5�6��^�#�7+K��]��<��J:,��f�t�+Km����������3�n:�)���n�3ffv��/vp,��N�%�"g\aۈ�����䢕�Vu�Ek�v�`ٸp�s��h�nNE�o�2��}�Ӹ��Ri���/m)^��&��]��]*z�c���7�>�Ez�k�0d�`��p<ˇ��1�ïJ ��XG�N3�p���>�1�ٜ�^;媥zجy��r�kdwi�C�@�����f¶KQ��i~B����l�^��da�����k�*���h=]v�Rw� ~���©/�Ay�ܛH<}?<!<�2f��
�P �³�C�vI�Is����`�	F��\$�@  ��[kuW���.v�l����	���â^	�ϊ����ޟ,P)�@��y�5oB�Zx����BSm5��8�̎խ[F�S�)�2	�񬈢n���X����sӡ�W��F��a����y�~�px�� �Y�ۤ!ϥ��BLD��S"g���E��+(&7J��T����F~���R�Ӌ����]��ج:l�+�����a���t�c����b�4Z���>NRl�|fG�lP��7'���D������o_<3t��?"
��8��G��h��"�D~r�p������KK�Jb|^l��I�����s 5I�F�bZ��[�Y6b��)*.�bv=�
)�#�%�<�@�US�E��d�sݽ�|���/�y|�v,&��p�L�8�a����d'�T��nE��T����M%��9|e7^��;���v�1?��R�XViZ��y�;'�d)�����z��I��fYP��)JV�]��1�m�3����#"�N5�2	��LR�<.���_�p��	�����y���Yޔ���?�z��~������2{��C�͐e7����b8|ޏ��/��!19��'k�T�����ˑ�2U*֢p�|�;f�����RU#R������#ir������9��'0�0'�&��%m��wD>=��y9e����G3���~�'�u��+�L��3gĵ�G\[,�Uێ��c���+��Y���_�e �5
�Qw�h#���=�/Ή6	caaI���L_�:)��v����
�� ƕ����u���uv�@�؝.;U0;�w1�ăw�Ǆ��E���_:�88�}O*�}���W)o��E�ݴI�HiY���k�m��S%X̔���ǃr�j6��v���w��+5�T�q/��O�1W������
�O�ռ M�(7�{q4 ?�2�)���(�?e�(��hBr���W�
�)�6�ĕ���'c<���2w���T�ŚZK���:�&x4��ܾ��������m�?�1����o�z֜Ҵ�C1�z0���0��w}D�$�����㝳�����#oJ0	��7KB��>Ȥ�a��'�Q�@���ɷ�w�_{�V�)���S�#M��h_����X�c�x�D�za}�"����SS�l76�; �;���˨�>��bp�n��rv���ƤM������Q���;�i��dc7��0E&X��{a������o�j]}�5��N���?*fd����H�`���_�[�����0��Tv9�[�qf,R*��q��r���^:�{ӷn�$��-�ldkD^Y[�SI�6�w���2�m��M�ñ�Koݟ�NF'�%�lU�
0'N��/�<�e�ǹL�LޒY3ba�P�B3k
��{e��+��=?=�%�;c�� ��X%m�ۛ�v�>�3	�Hg矖K����&������1��p)��K$>����R6�����k�����5.}�,T�����bO�o>Ü�Etf8�A���o[1S���)_ԯ�� cw���&��vم�<6H��ԋ��<3��<n
ftu^�$��(�V��JG(�.P+"w��a��g������1xF�	�ҩ����}U�9�����]�q?�2_k�&������l���e[&H�]���c��4�����U:0~���CBU�V�0����m9����R�����,�(>�ZL:� �l��&O˲(����'��VJj��tP5^���`S�uS�㴽\ijss���H���Ԃ�Ui��
E����ޞ��c��̆u�`Q/�ߵ��7��&��DDRc��@Z�¸��rM�c6�-� V=�P:m����|#�����Bȵ�g����L�d��@���y^} j�ܬ�%��P�q���uE���|��O�n#K;�	�"G������QΝYW;�/�2��%=|�%^�3qӶU�'J=�E�ya�ϻS\ �h�e�E��C�G�Q�_jE&��)�R��-��G��v��O[U��pf�5e1�����Vf�P�6�ά�ǲ&��̘���޵��q��#��b�ջ"|O��U�����(]�a�&n �u��]�>||dL���K$/��mE8Q�*��nO��ͯ�Hj�5<i���vL�k�{��q���?L���_��N��B	�L���B�Aʂ��r�2��@F-a!�E6;$���ø�ݎ���m��M@s��ȳ<'���b�ϝg���Evm���|�+�f;K�W������j
{:�,��Q�L�N �ٷ~�U2��g��+�V�F9玄��6B��V�����*���Aw�"h�8�v���l�C0�l�I�A!>V��ƙȺ�>��^g+����P�C��F�Nb:�=�8W�o#ϩ)!Q�T`,�(%E�{��nYA�Tƅ;&З���Ӌx�A2ਨ�1�P:���j�5v�f�.U&�e~�x9Gi����q��|�u1\���>�@D��U���'�@���N�C�� -
�"�[Ϟ�ol�P��moo�����mO��6n�m�.��Z�]��Lp�|[�1f�R�J��cofA㱲6��)��3��i�ݧ!��X��a���k1���	�}JIy�,��X~�K`ߪl�'A�b�%R����x�e���1g�ǎI��/��xe����|BP�����DRwd�qqOMÜ��@��-��σd���1$��2��cd���*�9�;6{�[~j�k��X�i�6����m���{
aOpM&ԩ:+=	G�7��7��D���b����hF����r�^��2�>"��}�����#� X�;��#x߂ u���!��T껩D<"i�����b�e������~���Y��7$}Xdg�ף&��Y
�UFQ�s��=�u�T|#/��B��)�o�^�����T:�X��b����i "�I��#�.��P�
p%w"�Ł�4Ȑh�� z�u���k��	/O>���H�A
/�~^a�����-]�P$b�4W!
i\nFʵR3�'���fz���S���oT�-�Y�|}�ƞ75.s���τ�����]	wU	�Q!��O)��) [��b�V�͛��п_?���N������(LiG-��E���Q֭�kA\�b?�ȝ���O�`xtg�YRV�Ն�i�ZR��e��S��bI�ZC�>"V}��K!��-�Vc����:狾*pR욍l�I]�&jzppC_+�e_�h�)"�H�>�*��x���Y/z$x���q����g����3�E���(��T���bB�v�`t��fb�l��Kċϻ������`N�_a�j�@�����̛�G�Y���j�l���蹍-X=���JgH�4����H�N�}9��	Պ/k�^"h�ksyM����q^��E�E�A1)��q���)�|#W�	�_�g~VR/�
�gu��c�5�	0�ʥ(a����n���|���a������]d0���#-�	��e�M@%(
ဂ��"�o0�ୃ�绦��Y5� Țc3�����v��#�?h��c&9�@�H͵��uN�����$�c��"�^�\8����C�3��O.a��2лc?X�h��\�y��sÙ�Ǔ�n�����λ����{�?�H�:D���3�{��Ø��)��IaX�N��)l�����K"��%"�V��p���D�n�C|6B�����̬Y
.F�����ٙj`l�-�ɛB/QH\���]�&WǓ�������gsv��þ�V[ERE5�_X����`���5^,}7��BIa��
+�<��:����Q�7sr%7��GGGY�*Ԯ���wT慑�¬>�}����6��� 3bD���94(.8���l��9�R���M�CFu��k��w�Q��K(D"a��۷o'gc$���6����&��[|�;z�!�=��t�^�9�^L��!"Jq���DFg�9��L�Z�|��xջ	ő��o?��[#��z+R���A����M�xEև�=�t��.j��b��F���9�
.-e@�"�	�ٛ�eb�-3~4�t�V�s�h��c�?���-
/h��%��)��i���F:�n	���E$���W@�E��s��C�w�s�����9g�}gޙ]��,7ãy���f&L��A����kGĂ����3�'��+
�����yg� m��sr/7V�D�l�4Qb�c��U	@t��zF�[f���c����5hv�IM����)ӑ*Y�.�#>�D+�m�՘$�2�l�Ҏf��A�E,��A7gH���Pவ4�D��T'������i��Q�HCs�J0��O�X�fQyQ_]@��tf҅��r�,��o#����Y/����KRBTVP� ��+����>��K~KȏwDMw54�C0.�M9H�5guH�vwI#�����)k��:&J��j;y�~w��8�H5�=�X�Ӓ3~�1~����y�7S��?��/+��w����>SIz��y��ja �jR�.�<>bHݜ� �pUI˿x���gƆ��� v�MNܟ�W�Z�Fr "�FM+U��(��SLh!OPŠ�z����6{��نIuȡ@fw�̫!b��������ʹe6n�+Ղ��3fهN1��d�¢p#�|+˹���30{Ek+��=sp���W#���ȃ��a9Qx{�K�N�P���C���e�E!M ��� �\(a�/t>�r�}�$9�������=ə�,�_E��ǜ�{M3%"�:���Rf�+I�@�`Bx��L��3�6W�1�����4d\�Ȭ� Y4�$w;���ndH��
����O��&�n�p��PV����H�����������a9"&�<��d�+X�2�,8(�j��v�C�}율����2�i��	�8�j�&S�Ɨ������Z�<�.�#@Qr.�'Ǣ+�o��^\�)_(�V�%�hk|��S\H��2�����/j�{xƊ�M6�坞Y�_�/i��)�6�e��B��n�����x}fA�ڄJ��0���Dkݷ�p?8����K�u ��\�O�z�w}"3y�J�o߆�+��|@�dHM)+)�Nb���i�9u��}�����#�#W�ؠ3�&�t�����r'��[���K��Fh�UQ�?�^���ktb���(�H�Te,��D��m�J�� B�T.�
�/�C�v\�	Dr=�8㣷�����Dg;�����]!grȕ���a�+�7b�<�[�(T�E���_��[�sF�Ѿ��Z΀���5w��7��%��)�l��t�.���&{��6/zOɄ�jQAi�֑5,�8A�E\ݬ�-�6掼��*��l��7%�Ć�"�� �V� +��)�N��5
2H�y_����SdDʆ}^�'�̷���/���~M�d�2�u�6��V�sC��ہݏ����$�7�~�����# c��\_f���m�@��o�~)��&)�A󈞩���y�����$4�6���~����/2&�cֹ7�䋉.��W���+@��j?�f��|VI�OJ�ǂTũ��Z���f�y��_�\]I �#/��˲9M�mA���E~����X��@閎��z^(}(&��_@�����F$�Nhc�m�n���^��$�8�e�/G�L\*��~��N0��bHyqG��a�`F�*�@1���*uq��#
����Z��nB�\A^�`�fL,]v�Kc@he�Z>R��������~:`��=2����=AC�������$�]����2!-���J�@?�l��C��� ���WS�2���qz�u�WOw����'$����Se�Lp�$�'��($H*)	��l=/f3���q��"�����C�qNe;;�oEƛ�A�䜌 u���'�3�����7��xH3].NR���g?]癘��1��&�FI����L����ֶ�D���b'�B����_L��[ٴ"(��B��g�y��q!W�d��FmP7L��N���U]OƷ�Y�I�._����F?����
Pͣ����Sh�2��I�A����*	-�*X�i���-��UZ�弩$\�rr��O���p�u(�,6�+9J#���o79�^��ї;���e�CIơ�� ��{�t��{#�K��#��ZZI077��;�wB�ƂA|ov0����N�gn�Ҷ)У����oo����Ɂ�n�����&�ם�0���G��U�kL�A��W�,�%��;�/s06L����,�����1,���EA^��+Y�4BZ���_�6��&V�Z������	��������F&���¸R�n	�zV1��"�y�o6��Q6��\��n���e_��#(5��
;����8�d7�9��/�:���2�>�å��c��r�!�r4���Ke��{#k����B�_�B��z����]8"}3*���u�6�qrds��9�b<�.=�|��0,|$�n-�q������)�ԓ_ �u=Yn�{�T��Ǳkal�|�kZn��'+h�=�5| �An0���>�2W����ι?֋���mꀷ�06l�?Pa�8D��5g�B�6:0)?U�Ƈ��״ߨ������W2�$�&��;C4f��(WC���v��@Xs�Z(��#�������k�*�Xvz���;(w�Q� �s5�f�cb���8�y�f�1�_��Ղ�z�@����uvfE�"�l��8��4� ��	#�k���h�\���}���"����ra���71G	�6�{h�C�D��ְ���'Ό�������@�ń�;��j��s���_E�4��:eW�xT��f�(�9>a&%����y*R�PH(v�Ib�(�����Z��,�x!��"����k{������k��/P ��k1��ۧo�.C�`��k�Ab�e�7o��J.��4^^1r-���>RA�[���aL��V��] H�_=�D�D)R(F6���1�N�k�ڭx���Ȗ���Q02�2���0yy;z�y��ѫ���	������ޮѬ��XQf�\�@Dƍ=�bf��P�������9�{
��+<����GpfM~e���O������J�QG�yfC�L��ۯs�)����ɝ���?Ycq�aw��� y�:��`��ʡ�O������I����~G1��&�a��G^10��f�"�)���?F���Y�B>���<K�=$��ch��x7o��}������زz�[4�8�[(|���7��Bt'$�~�y�dݔTj���m8C�5����9������J�v�R�{���� ��돘�z��Ik�.���K�2�G˺�[_-Y����ٟv*��\�Dys�-'�(V��w��".K�yR�������N�}�.��O��X�#���t�7KތxwcF���W�����M�����'���?=�n�S�(1*^���mSx��V����:��f��f�����AG��~�[�,��������E�z�]��14J��{��fѕE�	���N��.I���b�D���5��szzX����jzv� �eHC��@����-�w�,'���G<���r�_|g�<\o}�e_��h:r�g��� tkG737�{Ԇ&����=�f��H��786������`ڞ��iR��Gig�~�SB��/��h0D��悮��ݽ��c87c~���KU��f��x�K�(�$)ކ]+����e�ʩz?�,�B��!?�b�����������k��d=U0�h�6�G�&'&>"����A�ÔYN_��W=�
TU\�ּ�������sh��y}Ͱ=��͜?/�]�_����;d��N9��l&O=�� ���,�QF�@���e�(.m��Om��|~����a��
4δZ�c�׮Ť��qb7X�]b�FD�5�e!_��s�Ӊ��(��R�P�F
t��bi��=C(����~���G?#�M~�e��Z���\Bb ��QFQ4�������߇M<��6�\V[Foh�*0z���ՙ��͉Pr�2�F	�Z+��`%	x7�G�lK�--�:�����$�l7N�	�]��y	޸���m�]yxS�e�y��c*"�NN� ���`��,:h/�*�F�����.Z�?�)�����%�MK
:��^����aR��.�TA�"Bq���6��l��v,^P�ŉ�ר��xAw܇���DzX7�88�Ѣ��\"�q����ܶ�2'+�q�ܴ�����7�`p�7\�[:��J.��P	%��}���\˴�pR�\����y�O�x�zk@����=�A���;3��/�6?�5�rm�Ť	���1�m���0���7��\c��YZvm��vA%ȫ|��~sݜ�{<���f~0s�U���uW��q)��vsF�S',�rx�����5�`�ʗ�}&?����3S��zJF��r�c냐���.A��	S6Ipc�ɉ�߱f]p�P�.�����F��(��
�o��v:;�x�%�X�H��c�M%<9��?����n4�F��gXՉ
��tP�_�7C�e,*KA���үj�XބIp���)���F4htu�$��.&[�^��)��G�}�C��z��h/�����[���Bs��?�k�XI�u��#'���8�fi�c;�9�\�y����OT��$����b�?so��?���llN�7�O����]��X���E_ ���^dQ�!�g|zQ�� 6�{�+����_ߖ1�>�R�F.�ٴ/-�Fi9�4���9=h��l�";��mH���d�&�S�&
&t�����U�ܷ���|顓'Ev?Q��ʨ�X�1s��p=�������&���f��UC�V�T-���a��2/�{Nvޠ���eӟ1�E�zN�~>ex4*/�i�kQ)�Ġm���[�X��Ἱ��y��ML��;O�h�Wu��l���^/�(��Td�M�
T����+�������+�9{����F���x^�����n��8�1�Qhk@�؞�	&�"9��Ӥ[��t���TG��}����5�����b[��d@��ۈL�%@%���-Z�U��M�8ei�]�����򧀮^������'2Ü�?vK��P��cנ���7�����3o��Gñ~9MK�)�呻�E�@0�����aA%�����Q����m_T�����m�~g�>��311�Ľb�3v��3��q�)�����2x��$���O�ٕ�؞�pdH�n�����'EÌv�m,����<�!���kY�"�Jw�v^��=�Q<��e��/�4R�Ad�9���\�O/%��sZ�Yh@�:kr���	�H4��}x�2�VR3�����-�
�=
�C���\�a�z����k��o�y�Ttnk�[`Y;��kE��nE��&_����v����pb�q�0�ɵH>٘��}-A�\�����B)�9�Ҧ�Fo�;�}wG���p4.�L���e�w<>|V�B�4��z=`7��p����ڼ�޲GQTkhGD&��b����6�xeE��0�%9k�'Q����F�Ү-�r�"-y���=�vܡsrO���c�*�.1b$�bZ�Ȓ��j��tY�:��om0�1yg혡�����ֶ�D�tȕ'H�L)��ɖ�_!��_����g�:�/�ާ���
A�!B�;�\mg5�"���=�� ��/�����h�x$��z�j*�p꣸�;a�V@7-1@K~�m�	�	��b��X����O6+ݿ��n,�L�<�����������|�������?��� �Y��|?2WgER��1�����tX�@������
a�����b4��΂֯���H�je2��Aar���X0� ��3s�oR��_��
��D�Ѯ�O'>��7���#"�þ�D���2��`���ȫ�T�Z�QlݝbJv�ܰBϭ��d�v�JW�*�?,�Qȡ�����,�M��Z��	
��k���`����9bH�]��fz}�n�ǻ9@#�	/��U���/$�>+��}���1�)���9�=�u��=�%�m�`K��h���bɿFe�S0dEj�  ����[~���Y��r����j�kKĳ�nfP�jZ1���E3L��z��د�`A���Oۦ���0�s����C3z�Y�S�	uΛ��H����}�;6�Υ=���<�/y�-!�h�<Cj�^P�w/*�dw��1_KJJ�~�{{E���(�Y���1�'<<"�:�O<:KO����J F���\d�d�� s}�sO�+��C+���2�s>�Zy_띓��	*�2t�o���u�^�{|HL"D�;��f���{���❫+^�����wwbޫ��jϖ�ʶ7�i�7��7�^3�Y�=qaD���e��e�ma�w)΀޷��+��Q��ӫ��&��L�B�x�#��ee���j=�\��Pܒjt=ǰ�����Lm����Q�ʠ�O2E��$Kϴ����8:����/s��H�D��&>3'.OOУ��Y������m&�淝/O�}�`,��w���r��_���AUѿ�(e4�S�!LL��� L�B%�C�:Ǜ!1I���<�HN$p�����A5{T��/_���j�3�gr�n�	�
��|J���㾘S������x$�a6�i.����ԋI�ٚ�T�-¥w�ƌn쎯-OcBv*���(;L���7e��;ʵ�s�o(�X�4�����lֵ�m/����ߦ�nt�g�r�y��ҚqYS�o��l\��opݡ�{�;Q��*2�e��O^�@
�Z7st�f��ve�n�s4�`���;�+����*��J����a��\�K��w�Zh�Nk�iŲ����~��I`�r�3]6;ǔ���\GDN�2s}�6�`,��	y�aS����]�-Tf�U�Em	���RF�C��O
:~��a�N�TG��3�( %y�����}�����7<i����VvK+,l�^���o�͋ �������*A���J?�ǧ �V||�3]�[�����
#��C��,T����7�񦫲�S��ɣ��+��(�L�?(�ׄ�"멖3s'Nؑ��@(���Xj��@�H7�e��߿m�y��'�م���H��!D�=>MS(�F;���x�.$C\��P��;���T��Y���eqO�h&��D#���=֟�M���)J�ݰ�z#�a�n;�J&E�mU��11-R�$�X��1��7.�'�x��٤[��YR�Yj��/H-�=��+���+�?a���|��G�Ĉw�����K�?���"T�t�9o����)�ᬡ! c�N?����dnyA���V�_��ý�F���B,�2��׸Dn�y�wK?K=put��N��Ut<T���<�=��E>^�D���`�W����yG���Ug�z�ʩ�6(��F�F'$
7�>�Cл��Yg5!�bt6o�RPҗZ���ժ�O�r�����ͫs��q�N�B���t5���3B�Z���]��J_�!��R ��D�?�~���𗜜]ם�����:	��ej������G�m��!��7T�h�&�z��Ō�(�t�811�,1����Ṯ[T��\G��eex�c�4Y�7`��]�><���-��d�mu�Hk���S:n���~r�s�g%�4i��鼅E�4!�!Y�Jo�����w�����^���v��u����:�s'�8��|�e�|jI��������R�M$~�L��L�sk�P�#��j�G���0�~��Q]J��4ؔb&$Dft��oq��ܸ׺�|(��|�#���	�����Cʇv�Z_�Y�5�����l�����K�ρǸ�dv_5U����n�H���["#������5a��`�0*:(Ϣĕ����ו�X���$�$bk��h��(�ȑ��q%��L���^>��,�϶p�q->.4�:}(�a��;�w�d���(�kǳOK�_| ��i�)Ԙ���@F��F�MF��[�S� {Q��=�o��5���8^����m����8�Н�6����1����*/�_��YR�EzB]�ۓ�3<�$X�_�Ԗ2�D�Z�Y� M�Č�P��b�:�5B��Pٷ�g�)�Wʐ\�W��Vh�0�?@7��d��y�(3:�'��B����H����{�1QE`;Q�`� 0�>��N���W:�B�u訶Y�􎦽z[D�5/��#�5���	wzի��B�<U$�V�A��1�C�#T��,�}�j�=x*W�iy��w	��m���k����2����nJI�Π�}�0�r�MpgI��/7��!ܹ��tr�M9���4"o�yyI�%r�}Z���'3�I�������N���ļ��3����n����VL���8���19!�`��}B��S��jm��5���ଳ�,�"];f�n��&�t��d{CO�Q[$XX�j�F0��5�K���>��*}&g�)��݆;~�E�t�;C7�#\?�Pg���ڷ�n&]'��]�4�2�u�k���P��p�dX�P�WO�W����K�!_T�4'@�D%IZA#d����M/�S9���CE��_�����V̑��RsO��x��|��z�"�=<o�2�sr/*�;����wM�{(�����	��#%��-�~��>]ϫHuv?����$�ň��eP�>�1yfa�Ӛ���1ҷ���B��JJo�P!Uԏs�p1qE�r���w�Ȟ2�����A&��{z�_ua�5"}����H.�Bɜ6-��>�va���H��MZ���w_W�H���XD���,�~����~ 9�����X������t�9c���r)y����y�=����Uի��_X1����2=2�jO���q�Xi�w���~8D�ޭ=�in�akA���vbo��p�O-��(zn�	��"��nSK������׿�l��_�dq��߿K��j��Ve�J �fc��K�T�H����k���$�Q)\T!���L�����lԘ�+E�~�K3*��vJa�^%{1uk�]����m�w���c�e���ή�,֎�i
~>%d�;�)�\� ��8�p<�L�d�Z���W�Q0�����u(s��̈!�ً%'���A
�'�0����J�����EUx7 ���Ǎq=�ʺ��)�m�ȓ����"��ݴ�#G)�T!R�d�h{m=�Ht�,�kQ�TP���g����X�Ł��l��v��v��ϕ�@8��K��<��/;��Z�_�!%p�V�*�Ł���o���(ʸ�,M�F
S�5X��d�����ԣe��^Q
�
���T<�S��|� :�ҥ�f0sO+��a�l`�דgW�"�!g�R=��xT��8�дx�~�s[�����/���U��l�ԃ5��9�h���M�"%��*8�U������y=��J�*�FI��#�7��c�aJ�ѢG_��q�._��0��l�V.|Oq�'[N�H�e<�?V��wi�,K��D��=�@�&�O�]�jS9c**�\���wah5
﷗�xm���+hsc���c��xIQ�;�J�grO� �0�E+�ע�!� H�M�s�I�b�;�P��7)�Ze!���:����,8���"��
�"3��n�Pk�R�j 2�_cV ~�����C�O>���l�y����\�w����+�G�Ҵa� �"°"%�^c��D}Ao�,�Ot��K��5�����]kdp��kՌ�{;=�M��|�t���R
Α�c���i�D�Y�����9"zR�B2џ��D����ֲ�N9�$�c�8�Y+��8 S��..�g��%,�'3���1�_��Z������bԸdg����3�m�7EY7� �xZg�[
�+ӌ��5���-a�O�cL���*�}�������%�Ym`X}N��T*����=�ޛяN�H��n˽�.�;6�45-��aԉ��c�[��3�YcL�	u��u)+�ح��ִ[Ġj8R������Ӝ�s�FԇJJ���`�(�^i������m��y���ЮA�������܎C֏A?e�.���H+�A�I��7e�nFa2���u+gi��2c�㉄>%�o�cZV����c˃c)���M$mh/���p�b��Du�(�ǒ'H$�.8 u24*W�o�"K0���p�馔��xt���Ʀu�Kj��x�Ԃ������d��6&ЦA���⮫+���-�&�{_�������g!���� ���c�|M����"�(c��ġ�@*bk�ږ��Xɯ��(�j��[ًےx���iAߝ���F�s�Q��D�7�Dہ�L����ڟ�T3�"e�o�(��8�y�"v����ck �L�b9%��\�ۇ�{��S��+�Pd _4�N_�兄`�'D*U�.�x|�6xY�@ߖ�c��ة���U����=�
��^{��T�Y(N�ͫ���
�a����v���K���[�M�Z��j��ӣ��tX�J�ѫ$Ký�j���
�0hs��~���zu[��V���r�	�;����XSL�1�Eu���~�WM�%	��ZF1����p$5g�����9��__dU^��̬�ڍԒ���eyd�R��ɖL��Q��^�o�c��_�\J��6+��c ��lŉ�?�jW�%0��gh��>N��&�W�ࠈ=�������L ��È���\�WnF����$I�@"m�W��߫��3�+�	�TD�����G�	J�qնծ����@�g�Cv�3��bu�(h��)"ws���cH����Uc��_o2pglOE���/����2��Y0c��gC
q�5�m��e�[�nrk�orY�4��s��~4�A���3	�l��y< Q�x���#ŉ�Î�z_.���3�d�� �ײmـ�`��ӝ�J\|�,�ֻ������k��^I�"i�O�ė����	Y+C���v�. |�K(���H:a񛯆"�;Ih��s����%k�ؓv3��}���1� �AcvU�b��(ɿ��ըs־��%[`!u<�Hc�ೞ��Ć�egzZ|�{��&#��/Mk��A���lQ̀�bXO�v���L(�.�J�+70���������7���x��
�?�}.�1o���CuF_/{������E��_P?�@�ے�ë���#�O\�U�
U)�F?W�%Y����_z�~��!L其�t{(B3����}]Κ��ЏK.��^����ci<~��?$�&Y	����!��d��^@]�c?e���\�@���98��fZ%|��C�1Ek"d\����]�����%�M�[Zh/2ܙ��Ԗ����������@�e���������/��N�W�����R�m�߰�?cxz�^���}es��-�p�ΝM��ۼ���o�K9�.�����S��x�޴�}q�r��[�_Fywr�EUTZَ�d3*i�;��jE�� ��ʓ�v=�bv�uf�����;>=�s@$��we�_�<�iK߱��--�O8"~/�wn�u�d��o�u�`ߓ���� ��������Kj�e@��p�u��v��GV�.Y��}�L����Q˝m883��aF�xnX_eP�@�ѡ(鼠�Vr^_�t�C!jC�����WB�����A\}��ݷD��=?�Y���Z���g���h�b�C�	�|�67o��3nd(/�g�jC�3�{���7�k+��Iy^�o�0����T2C�@��(s4^���~��+�ִ.8� ��RQ�5�ľ@��,>�i�A5�p�7���8_/7���W�׵5�@� $��O����VTI��O��P���N�1��F�(P�v��z�����Hxo��ɷ$r����k-K��V��8/��F�#8(����|��(��qO��;����p���1״מ�sA�4�Mg���J�.s�@H��.V����b;ja�Mˇ���;�w~W�)ez�GO�
��>���ۈ��
0L��D	���"�j�q#@WP��z�ꑾ<�7�޸���|��j�F=���16H�@<w�"��@ø�43|��ˌ�W�LŔI���q�|����"!���Z;�z��tr��� ��b/f�V��j�g߶].֪�D�Lop�vTr����ˮY�E�=&���������2�s�q�l
���f˕-��Hv ��ijW8��b���,�x��vi{�s� Y^��O���=6���*�r�����i�p��0%3�r84vD�H�ֆ�֥kv�S� l�j����+��`����勬�f�f�����G�~�x�Q���+���6
��)*�{�`��.���J  �=��ktD���a��Xc麉��|�ڻט(ƶ]hP��5w�&��͋0gd;[�W���d�q��l?y]��,:FԠv�F�BpG=�����b̌��L��R�Z^I޽ǉb�<eC7�<0�1�����9�W/0��T������=�&�UT�-Q�W��Py��6�O�XT����1}�>^�[�wz���}���G	��!A��]r���K��D�Jg�Ϋ�Mu�ԛ��{����L""��,� [����TT_��ؕ��~ֿ5�;M�|s����׆��bq��;A�撋�)�����\���<G��$~0*d�럨4�[�X4��p����+|��C����E|�%�G��/�>�g���
��?ނ�|b���Z7��������#QלP���޴�O�	��YK�gu�����r���B-���� aU����-G�/[��=6���#�F��z�~��ϰ��B�J�5�F0,t����� d��V����[����fY�[u#�P�t�Ǩ��n/����*o��`o�
 j�=������v�%�E�T)�_l�9��Z��{,~��{���	H�Y-uh���`��I٪���t �[d�����*�qs���b�4��Dc'�A�~�`ƀPݔ�������)�^$����W��G�j3����&;ʹ��8�P�r��J�|�'�F2>���_D��m�61�S�)��ЃKɆ�t�x�"�k�.ėyie��B"���h��W��y)��vz��[[���$ia�*j�˯ƹ�3bozɾ�xz�E�։�bmc�lIS�6���=��Q�Y��{qm��^�WY9���(���s��h��=�2��� T�I�%����??�<��3�Wvm���>�o���f�:�<���cU�����>�˥��S��𐕱�S
�p+�,�j.SYy��>���|�Z��U���Qc�P�rs:(�������l;�тC]���\�f0�U���c�-"��Q�<��E1&;�ϩDG^'�/S@����z;��.���C�gg>������4��א]���*~s[-y~[N���Ɖ7*+�{1k��W5C� ��Sr\��\�~8w��#=�,?ҙȫ����	��1�zX����LiD��.�ı
X�$n��@W�[Et~��C�����o��B��Gp�:�ΏE�e�TYn����N�'k�}�4�Z^���g��!��$�ArӘt��3��gJ�7k���������m.��oG5��CIFz׍w���o����'��;�Q�lT���jL���u��;�͵5�Ti(֑���Ҿ������2d9��{=�Nn������� RP嬮�����`6�&�ƮS
B�zC�$f��~�̆^�z7�����>�_�rbCP�l�2U��)`����I���� �F���x�]�j=C��1wgU AoY�s���+�{��׾���W���;"^�Y�� �a�����������<n�}�IM]��?Ytx2���v�B�c�s�v����)(��Is]�zO�q_���Sb��* $���Ivy���X�S��|�3�F4�{¼jHۧ|䕅�i�<��/U��X��������+P��s <T�\y�5�w�+u\�n���2Ĵ��)�	�h˔T��A+�"n�ڒ&�n���>GF�yԦ��={(e�8F���Dh֨�MzM}�Zi������VJѬ����Q�`��F|?)�����N?nfn��|�2P�j?���3��n9wqe�I�_��m��_,8���fz�Wĭ����4��K�6�tw�c�PG��6~�����3\P@��Bs���k��p(��r�\�+���!�)�>�.��/T�5M<hY�YhيG�H����ǣ�c1��X^��Ջ�a#�%���H�o��˞@���	:�T�kii�`#'[��j����bt��]% ��99y@rh���(��JΦ��m�%�,�k���^������K&G�g|��G�bX�I��ϡ���U��ˇ�ˇ%WZ`�����!��z`{�d*l�7����Ǧ��|4�8���ן�;��`��g9��@,�j�Mݶ�X�sC�f��;S�5�> �Q����̈�t����:���wDc�tCʃ&�����4±�ũ\x@�?ob$N?�#|�r�����GMR�{8}�x��p�^ٍ�3�1����<�r	�a�9�q1k��7��X��P�k��mc��rw���#�]�9\�٤~�$ߐ5��0�nڑ�m���PyX��M6��&߭֜���?�	�?�,ۍ�Q{�	\��3�aF&�*�{A?�ݧeK�LJv(��������"{��}95ߡ=X����j����N���m�eh����14���}�l�9�ƈT_)0���z#5*?N�$UG��K�AO?�n���������?^"���ڵ�ҏ��Uv���k����5fxC��y���'���Ub/��i	܉�
vnH�+í`>�%���UFa�l��V�CŪ��
/ù��S�d7]�|-:ߒj8O+jA�&�	����;E�PW[ #&D��D���.�?�uTg>�zB�d��ژEJ����9��u.�-;������Q��\��8��X��L��z�C.�C���3`��q�Y���8�~٘�⹊!@zt��6H7H�ҩ���`"(�&E �~v0��x�Oe?R(KH�U�T����^��h�����>1�F�!�m��(\��k?���� S��3����-p����KJR���k�3*g��X����]`f��۬�e�'~��򏍣�Q'"���iP�g�L|��[��7s �Y�Y��@#\�]1����:�l_t%�״�Щ����`����Ff�{�R�(���F�c�P�{�p�W�(w���AZ���A���>��<n�׺�W\�&:��/�gT�/�t�)�ZCʡ��Ϟ��i�9��Al�	�Zp-����=W��n�rxe)�"0����З��FIA�梯�'{��;�|��B�츴b�Ol�X&�+7�s���J!D�}�ϓ���Y͵;�^7eo8�����a:�O�:sJ���d|�ԈŽm�\ߤ��>d�ES���L�_����n��U�^�뜦ӀNV�����u/�'�b��Ь�	[=��~�L>^���%O�����۰�wQ`�H���R�����x~��M�����#
ҫdօ4�(���nX3�A���׻u< 8A��R���砂�x0f.r݆���*�4_��m�ܻ�e}��A������j�Y�G�}4���]*���?\�5W��h��!�)��%[����sU���{Y������)��g�"�F�R��K�;��0NJ^���2� �l�q�\s��d��Fe�@{�UC�Z��m�-$��;Ə�����R���8�,H)�7��?a���A?�'[�`��	��{�!��G=Q�w��F��~��bXo��@ǫ ��+�ꈟ������B��t�-��9�������a()��"0P��[���*����Җk��/F	v>��N���7]Kαi��������Q��a70�f��C�q�<�s�&_���Z���yd3�kr$��3/8�?��v�Q��A��Al�}���)���<��NY,{H���k�'pA�!�Q�%/5�X�#`��G�C�i/[�d�R͞�Y_�ʭW�a	���J��WF^�[˥�6��E�r5���x����Ƹ��n�xW��dSJ-�e�`��m}\�l2F~{�c��c��q$��&~)�����q�f�ؐӗg͒؀վR�n�~5�7��E�P&������A������զ}�a���w}Ҩv�
��D�S�)o��kq��G�V���X���"%яz�������^��Iz��,6�ACz������,m�D�\:����RY<0Oc�Y����⫝��G�`�� ����O���՗��Fz~)	<~'���>�J�6W(Az��f�룩ʛ7����eUد�w�����;�HiHn�d�� ��e;Sٖ�c��'������� X���WcQ������D�]K9��ܙ��J_&�|J'��;%�)�͖� ]�C��+c2K�m/�!V���Y���O	�U8�q~!q���EJ�e!�C�֫��k^:b�V�F����PNS�A��Q�%"�?S��y�ڞ6�G�,�;�	�4��W�ɯ���0ea�﹛1��e�77 ��.�B�6�~�!�܄L�#���e���K%�\����}ۻ����>Z��IS � ���﫨���}��4.��١K�y�CT�H���M��w	�?�y~J��R���=�Z�I�[.�/z����k�}�>
��!-�nt��! ")-L�;�I��"�I�%%G#�!"�����}��cǳ羯�:��y?<�[HX�~��9���Y�>�pJ�J��;]�������f	�3�?��JN����H����Fݨ�?��<S���Ӣ�[���"1�m�vt����S�A��)Ż�"2�0_i��,)���k�p�Pki�df� ���i��?���Pý���x�d�v���!��E%��:�M-����jr���g�G�I����cuA��è˿�K��ǉ�`Vv]��C{��\W��/�T��7���dKw=s��ڼz����^t��"�� ��f�M�/YvxY�Q1��f[5S	98.��8�����9r���"�b";"j��^Z���_˩y�v��g.N<����s���T�f/�_�'��A@Y�leЭ�Qʯ�Z��Lϴ���B�|Z�U%{�ש�|�j�cZ��+��]P�%��k٘{Q�9�?� ྸ_��IZh��\�u�����c�tb#D-L_�ɈVs�˨=��y�]~+إ�]MZ öH��}ҁ�:����/˴+�6M�c�?|�trOᶀj�
"b���|)Ch��0�S��ׁ��H]�0M�]췝�ZǇ-�MGrM8�!A��~����⻌Od���T�֢W���g�֥�;����%���]�iR�)���!�O����p½��)��fwj:(l���l{���8�����Y�W�v�6�} ��{�pj�Qr�U�k90o���H���:���\��_�z��������?1�������$^�L�O�!{�褻������o�MNv��A/�;�������M�(�+�!f�\wsb�~����A���"0�R��-�f��ӵ�,�i���J�.6�菶�2t?�,�#�U�Z̸Z:�c��i�w�#�hYfbӤ��5t{h!Z��d�ǻ��#��s�G?N�9��e�"/�d�Զ"��0�t�s�u��Ɛ�'�a(����5DH	�}kw�g�L`x�gW��]�ER36RLYOk�m�j7}�'ǗG1�|hc�B��1	>����"K��Hd��[�w�}�ޮCZ��X�� Y���c��Vo�TԸv�_��0!��t)�u�@]Ig�{��}�^{�ij����5�t�U��0C�]O{��1k [���u�Л����)c'������@EB�{'(.�Q/1��v�P� d��t8�L&���&��NQ�7˃J��>%�{������ޛ�`�pi��r����͑�� J��}W�
�U:���MU0.'S�;�}��S��Ƕ�����!8㨕.��%�Y�F�97(*��R:[t)@Z[���ϰ���Ի� WryBK��ꥁEe4P��K!�0=�3�ӹ��t}�E��#4��xq����� ��&��kC߄!�YG��
W��c��I6��t	��8��4�'&*�M�+���*{�|8/��Mփ����L����2M�V�4e���}��ȸ��l��{��Ő�@F�	sW��uE�%��hTu����lC�Q�-2��+y g�no��Ӏ�piUC���T���=)��t/5dyp�z{G1�@�~�	���N@{�ˣb0UM����f�+�q�!9�#B�l��{�$�DF{��wX�ӻ�3%���Ƀ��v���wm��Wy�;~G��Fvv�'�R�G�~v���>���T&���9Ȥmͺqx/�L�8�A�����?�V�jb�CD�^����_胄�o�tFP������A�<fP�@|�����SQ���/�M�c"H������a8�]	뜶>��UK�u2��w���}5�C��E�����鋞Ö4hhr���|�Z���߶wY�${��W��}����z��d����`��l�#P�듫�wq#R����]����ZOŸ��H�9EG�����$;B�t��n[�p�p��t�5h�h����E�oX��b��aVt�8��6d��iM^{]+��w&ٮ%����QݱX�V�yw���"4��R�jc�n���{��g����@0q�����,���Ӽ�y1����cvrRM0>i��#MgD�k�^FK��ABoM?TRq*�3��=�o�����Z���	x�K�����	��i`���
 �ϝe�ʐ�NU68���-*�N��H����Y�S�x�B�>az�*%���!��B�8-��\���%�[����(��;��QCư���l�I�b��u������|�����ܵ�~E�g`����d',>Fމd�����L���c4���pG�3.��'��V`F4��>��"��I»(W1C�
�4��Kr�z�ۋ���[�2L"�K`~N��Y��N7�f&a?Vb{��t��D�:�_�Z!W�R��R��c���������`%C%���1:�&�(�{�4�������K�f���fO�I�����P���q1N�\����*�'.*���d̜H<h��賓����A�k��4�!��)eGH���3a��7�RzP��d� ÀÏ������=d����#Ⱦ��߸Nԗr-�a���vK����e�@8ϖ�Za�����S��΍�A\����̝ͯ��J_�o������u>�,
9h����x!to�Nز ʃ�ܶ��xL\�u��㏌]h�$���>�iw��l6j@���^3�F�Co{W�� Đ�˒b����B��H�������8�/�6��3��\�ӈ������h@���q��4�A*��^D&r$/t'&eF��A��?%�:m��<��/ւ?�4U�:8ΰ�զ/� @?�ׂe��oVx��Ty2_?�r�w�bm���>8;8CI̾著9T�ja��������A7��V.�YN�x����HZ���+�@���Q�����1�ek�>��Ji���!�o|�d��~~��=v��[P�! 'jR�	c �ކ�ZT<E�'��a���gX�Dߴ���s�; Pm�̮��5����2�AE�!X����	 .E
����OsR�=[��i�fLV�a��,�@q5�����ۻǆ82�U��v��f'�g1u]�%�<Q�@�_��0��Q'�}���N�ÿ�O��i��m}�)X�װ*�kcrG �L���kme䧘q�}�����ZC�'��ҏ*�������d��� ����ܯ�+)(�_I�Q!����< P�fK�oÚ���|�%�H;�d ����P���Y��*�A��O-Á���B�����YoN'����7�I�����`JHCK��i{�SE�=�� ���6E�%zkK]Ʃug����>%���I�1�#�L��`�`�A�u�q�^��TX���0\���_p^����in�#�7���P�Pt���0�Ye��z�f�}v|K��q�� �=�&h���B��Ek�����b��iP�#t�f����z���0�Z��`n�\p�����=Q7k&�@ɀ�H�W'.T3���G6�z	މ����*���Nx��ƌ^�Q��r����Y�����[�?�w��nQ^@5�q�$ɼh�����ޞ�W��0��q�yFL`�~�/�I(�]���Ӹ	�g,���������	u�b�y�mSX����y���6�b��>i��.Gl3e��ܯtK��/���&{�	���T���Vf8���Ggd��4k�Un�FO�{�>|���֞t���UB�O B?0ؼA?���Z�I�73&r��@ zIƥ]l��N� �rH�z_�z�b���r�v�I�U��8=�l�q��[,!������Y����������G�qh�me���~Xi�^"���Mm�#�2�8{t�MK�xX�>@�B����%�h��QxXm�!ks��3x7k�w�ysaō9ұ6��^�Ȼ�"�.h���]9���)�#x�߆4���7Yk�]�SS/=6�����cJ����-�}{�o7�3�J��������|�4�}Oe�d�"*Z�PO#w�����%�S�^g�yOᝬ����?�0s$@ X�rs־�s�F���6��  >5b�S����b�6^`���_����w�b���2����o�`�^ �NĆ����5E8��=�(ul�.���q��^h=*��~�]�W9l�T�#Nc�����ɼo��O����r���=��/>tU�b�mԉ� 2<.�r�&��'D�b�g�j*��l��ǔ�َ'�&��`�C��i]/�� ��ΰ�y���}�����E��R��e1�C0M&�"hn�:��8�65���<<��ڼ���>Gƌ��dأ����Xu�Nǭ���Ǆ��w�m��.�8�0L��<��0y���=Ql�Ł[���r(��Y�������Ц����#=�!@s��aދ{�+��G$��e�a��Uw`�vV4h���伃���t�<8В)H{6x���G�6�2�LД�����P�q9/���5�Y?R�g���!�iPT]��E��I�8_-L�A<f̡
:�j��t���`��ih�����Қ�>�%_����Q�C�~st����*��r�^��8��Y�U~rJʍ8���=�q����S��l�������9K���F����'�f�b��g�5+�0�)�4O��;�ז����i�����/�h\d��{B�}�)�lTI����$(��u/��f��m��zG�~�����[oW�)g�דl3�G�*:���B��w��C�&��ǿ��J~�t�&�נ�-����ǲ9b�i��`ߋf�t�����A���l��Kx��o۔�j��8����%�DtW����W��i�xN�O�F=����[ݒ���.�P�����|}k��w���l��:7`��_�u�~"��S��o@�pd���Ӭ��|���{,db�P}��q�5Y_��Q1GJr[�Qv�o�S���6�z�co!`�-��S�_����y��W�q�TRіFEz&п�_~�*��=�q�S$(�����F%q����i>�$�nSo���U"����ԅ�ӓ���j���_�Z��`����`h_cMP،#�B����g��&1��\b�*��b���ګ���?p��Vx�fS'�o��3sK��t��������;}�%�^�q��tlh ����o!%]⚢�ŀcM{*c�D���)�'��5��X��̶�^"~'�&q`	�*^��=EL�
�=��PC퉺��#�Ϻ*7�2�N��-��)�٣I�apW�lR}QiC�5:92��.�`���iȝδ��J�q~�=��4���r>�U�{���
j�z�%~��E\��x�?|�c�ض�;�@���^W���(����{"u �v��}���à��趖�r̕�H�.��Qs_��ҹL=�	姃��{$l��;)�����L�X֦�>�o|�"�|L֪�Z�4;89�\�~
]�	u���耸q���e�����foJ�������M���ܘR�YOM��kbʇ77��}�J>��K/�2HYr1�Y�w�����l}l�#�R+��?[���Sƹ	�w �p���$��y����Ð��L����h?��:ǹ����V�)&����|8!�)Y���
�U+ij!����Q�������N̐�.2�1�Z�_~U���Y�6Z���?~Q.r
F�a�]�v��+i�W�"u�ߦ���W#��؟k_�@[WDq��cS��m��i^�{�ZI��W�z��ж��I��+��{�^�U�dQ��徧J6s���gk"��F��3	�3�n9Әz��{R�g��{S�i^�Ⱦ�F�V�tn��f�}mq�UR.�;mX}���������z������C��X��4*��|���V���>�wD֓�i}8id���?�$A'�)��:�x)���>;�nE�d���%�뷖��`��x���wQ�C�4�&�쌎��#Ø!�1��tE++]W.9��DU{���P�/x}���ϼ֬�����˸��H��z� ��4��c�{݃�3t����h5u[���ڔ�&X$h���A��c�+ߩ?�����_�J�.�� h{��`��H6�����.�7��Sr����헥w���k�&N�D�?�LE��^QN���%r��:����ȝ�&���R�֗u����M
"������ꇢj.��G��)����T±೏���Cy��m5�B���Qa���:-��9�}���9��������뮮:��R���aIES;��nK�ܓCn�:Ed�����ɾ�2c�����Y��B-Ʀn��2��w�)ݟ���ѕ��M�6~�g��Y6F��L)����E\�AۗW'����3�LnB�C[��bU�y��ؚ
�y�����G�9Q�S�B�WL_��5����.zD��DΠ�p��zl8��m�/��$�rA���gܹ����_=`�h�b|����� �oPP����6�<r�DP͹����?T�W&���jH6E��;`G�Ư M�N��?4F
e��I���e��qy��7�Z��y��#?�fZ:�U��/6�
T��TpԿΐ�\A��Η����]eo9����C�$.)\.ݷnO�sG_�	�mՇ�:���:S^���1�q�2��u?5����~��:x�Q�!� q�k҈�%�mk���f�9�ϱ�*��:#��T�bܨ�����圫t>V�/T-yNM�/����H��ɬ�r�Կ?��<�`�wD���ɜ�eV8��p	"��&#9�,�DmF?��o��_�S����~�&��{����~1Z�_�}�ܩ���*��}e:�]q�$\&�(�#PL�ɶk�9M��{@7u���a��x� �7�M�p�#���0�bD�^�s�x�
U5�����u{�m�^⹚w�����~����S� ��;=�m������d�ZN��=V䗽�����F�X'�D^���jg[�l�9�:��=�1�����[�#CL{E��Ycc4�a�Y��Ie�����=�V���BڢKgМm�罖�kN������T��S���Ɗ�}�PO)=T��I��:������b�5�ᴕ���8Z��MDҋ���tO;���`�hV���3n!�>m>�ە�,��>��C���� x��av�*K��-�+�|a�u��ao�k/�V��2t��7=��t�U����o���""ӗ_�ˀ���_�گ�� o�]�� ǋB���V����B�0�굷>�Lؤ���;�:k킲`ǭxTѠ$[�%1�<1��t폚�0�^,�0.YԪ��~��jZ�LCvk�=�n�5^�J	�'��X�"N{c�Q�W�W݇����A\ ��7�iK27	9#|�&>
>�ݏj��Ƒ8i�&f�?�YP��r��#��N�VX��^�&����w�fث��ҏ���p��,4믋����������J@��l|`�:�5��y�!/U!c��j���%��y���%r� �OV��{�'팬���5zy�����|ق6�/���Xf��t)֠<ogAN�g��������"�ǲ�rBA�BĘ��E�V��5:P`�@�A���%�(Ǽ�;��'+�ɦk=Z��A�fVղ׃�]�AH����i���z�$�(�V4n�ߠ���r�*�It�9��,ҏ�x�`�`a�<q��.D�NQ�C��G
��Z���vV�foV���X��ڂ8����|��*j���N�����e��!g�4\�8Ch<AZR+>�^��&��/������i0)"E����8`1`M��rn��v��J6AQgT
 hk�)J>�ͽ��`��֊��]��½��V��|]�;�ꌲ⃭��*[N���R'���
ߛ�\���x�oe�~d�tK���� ���_hg�<��ߓ�����:�]w��uti��|��N��
�*I������&���.�V+���v�d��h���Ec�ZE�Q��Gà֐���i����\�����`ﺐ$]��k�ue� Cb���7��_
�$~ʡ!��"t�.��#�N�0�q�;�m��O�;6"dOZ�ź��m���F�;��N?���\$�M��*.=��b���"��	��A�p�,�0�E�������hQ����03��ӇT��L��
	��S��{�䙞�\~g��M^�����*G��|}i�j�5v_�34[���s3�rxk�`��}��)����bO�q������!�$�Dq�����zh��:ٯ��{�V��X"�N[~�y�N�j�O�~�[��r�o��31y[��R�ժ��Ѓ��E\�i�~�����*�5���a���1���������Uٴן���{��(m=��T�Ix8�p3��Ol�Br �(R�zشN{�>Y�7 ��-#�K��j��G�1کI���~��YO���X�;�Ә�N���m�nI�*Q�//W>�_6�|�Z���&�*`��0�[�~jUA5���
e5沇ݞH�V�8D�Y#��y�;�!@�~�`1��#<[�B~��a�޾Q�vi����w�!�,�6 {Y gߩ ȼR�|�8�g�%��/�|�Yq�3h���#�Ѿά����!��t��]�j�Ȓd����X�(:re)o��j���	C��oq0��<	�����#�M$�q�m�륜Z�@����=���w�B��FMrR��Oߟ��aoY��ԍ.4����5\���-��I��+�
�~��+��vivaQ�x,c���9�TJn�r����e�׃���,�!&��Ǩ_r�۠K�+�79�.R��E[��7<��x�D묳�-w�B�=�g{
q������<XE:X}�b�������"�Ǆ�s���s
�9�l�±P�a�*~/�o���;3XS�J�<B��L�Ej'\~��|�����K!L_M����)���_�Zn�E������3�h���Q�O�F�������ʝ�L�2����@�$E�n�?"Q�o��Œ�_u-���]cSW�<8��Y������`N�C��{Q>� ���S��>�����x��Z����+����v��T����妊�8Ŝ�o֒�Re�*�<�f���
ۯR8�~����![�^}y�pr��\�x$A*~�c~�ɷ/���|2��YC�&)�*$���-�`����3^R9�g�TH�n�e��`.�V���7oϭn��b/h�Q�	[�L��@
L�x���u�m�{w�G��c�7���lD�~H�d�6���aJ�ҫu0��z�mC���R�*b3�u��7���1����%�wcH��ǹڼ�w`W��d�m�Q���5B��)�Zz�WXLｼ=��g�z@���7�z03�):���Ĩ�m��'�h\�0�{K?��<��	��ZLz�������e1���	Zy(7$��-���^Y�\v�J�w���%7��T����ΰ}^Őb�P:p�'�����i<�G	�~$;PQ�W<h�ڢ/B_a�'4�
�t�����84��4��WOnA#�F0��h�J�ՙ-t��)���[�<�z���t���I��**��MQ�O����}�� `�G������+����4�U���Q�<¾j��!��S����:��C�V��U�"
�c9�ട����vr��*���n*#O:Wk�iKc�$-�X��� �t:c��:�0�(�i�TIG4��ݕ��~e{E���lr�t= Z~�Buj
�F��=y �@�f�I� {��,�\`ۚ$
����w{��g�qt*��\,S^b�t�������DҪ�1�� c�x����;�㠟L	����]><��#È��ަ�������4�9fS���" �5�o��h���HCj#�g1QD��'�����9&�e_G蒖Z�4;C
ʯ�Buɐ��-{ �*��g�s����R_n�&�~��C����()��u.T��d�g�}�`0�N����*��'D���6��펽�P�P�����%+#��������Ӊ��%D��ӥ\����ߘ��,�����֡�>{�&�Oo�ђ�id��<6|kK �#�$(��Q�
�`mW�{ҭ��G���@�D���}N_&�r���	`����M=��bFr�����¿�}[�����R8�����mMݛHA��I�J�H�ߤ�4:h�kiAg�k�d�����wna�C�F�i���ZzQ��N�w����§!Y0r�=k�9Z[;��Ym�)��������PN��(�2�=XOL�}}��e�gf�����nI�Ҍ'R:E�+l��b�U��'��D�l4��y�L���1i����30�#O�'��KE &D�ت{��b$�`�1V�	����B���E�D�o�+��ʮ'�]�G"O�K��������@Wm��������<��+\e M��v�E�$�E�0�%�5����s]D6*� ̛F�� iꍠ9��'����k�P�ӭq������@}��X��"z�����j�.�df����Ӎ��1I����e��s>!m��c͜�=�i� f۾\;�@�1Ko?�� `�]N�N�u��]��?R�s
��7g{�ߗx��0��+F�ú=�~�o�{v�y=�Ng�'ug�Gۻ���A׿�p\M���1'ܓ�p0�Po�CB�`f+L7#��@~�"���;�g���{��\�������I�����>{H4 ݭ�_��p��U��P��`J�K��F��P���Lqg6�Z�9vXR�֤�>v(hz�8����.T��Օ�������	����0��\Ė���y���浈�|�LN�>�M+tM*��|�s�L]�J�y���Nѡ�&
2
4w�;��3��-M2�C����|�>�c|���IGQݴ`��o�
�d����(���X	�Ꞩ[�<�b8&�|b�4�R?�+�W�~���C��
�Cw�Oi�a�œX9��e����	���h���t�߻�`&q*�}���o�:z�Ӿ�A��;��\�N��5�'dY�0�-B����q���ɔ���L�$�'����xr1?vY��O�'�l9#���w�&r�i����rf��?�H��.��H�O�3'N����bbPs�v���20P���ğ�+.���d�!�'*�5���1)��>��t���p;2$���7��p3�E>��e:z� �+'r�-�q!�.��� ��#�j�'����m���T��@1G����к����[�4�-)��17$�o�V���9����Z�|�����}�������!к��6�������P���-��Fz�m��m���=�e�����p�(a��gK�.�;O��$4I��wA��(I���E���?Ɖ	F�eE�'������7C���V-jL��n��x�+��ܭ���,�L^��ǲ���N��Ri8�d�O�L�E�E�,��(���IWr����i�ʌ�j�J;�(���~�B�GW�ӆ��c������%U�(�ﺾ�: <��X��#C3�����iE�ZG懽��xߦĔF���@�\(������3F-.�A$�J�PgMڹ`����,��E<�7�,5�:��V���0&W�k��G�Q�30����.w[D���5UQ��!����xl3�������g�+?���܋�R�?Z�F;��~K��uv(R�v��a�����A��ˋ6���D;����PxF�UXJ�pd����<u�{WjC����_t�t���|�KP ;��v!#�Q�����"���AY�fo���C�&in�52ma6�aU����)X�E��j]���
�|&��\��,Lf�l9��0+� �����}�z���%eӰ��k��}	x5T��,���ùeUz7�iԜ��ɥ�#�뙚�j�M�ɒ����@�Q�t�.��."�^S��/ʣ�*�qU:Iq�j��O=`���x�@��﹮�mĉ�x�7Sp	��ˣ6���sPf��BIs��|�l��y>Ea��:�|��ô`� �1ٓWi�n�����n�z��0��f63�rjaZ���Ov��ܗ��0�I�IB�4T��V�{���,[��S��|���]��I�}2�y{x��\���Ent	�+˵RGW�����9���)�Iא*�@�ʬ�h�
����'r���brMx󈟷&�4�b�QtA�|j���r���1B��R�P(��t��3T�]�#��K	=���,6�{5qC��g��##�\Ä	���D���f`8���h����B���4���P;6)�|��7*UK��]6<N\�8v& .�=�iJ�hgc��Έ�?��ސ�ؗV��W憝�[�߽ʢ}2�FC��.�t*�{�!'����;�8��ʡ ������?|���a��P�'�G`�V�~����i��	H�o5^�rm�����O��ӳ:�5J/�]����'�-����#�Y�G�9�=�>��3�#z<����f��������5~�#q���6���vc���uN��%��q�K��Vu��"�BpF��a1`�2�T��A����� �l����Q_|��~�u��L��������n2Ʋ��!�8x���H�XT�Nw�dŊ�K��1��^ʿ�5�e�S��޲$T��r����즅Ii֦�<�ڈ���@���~�G���>�HzQ)�-f�����AP��`r�7B�-ƒV І��^�))�`L��?��Z���A'�����sQ���RD�fP~��*��1�;l���ſ������YG����U~��Z���D�#��oߩ⣘���}����s�����S�*�k� +5����Ī˺:H�TH�2�?}�8��1�P���3(HC𨰅SI�i�,��H�Wp���S��I���1Zpbx�Ru�:�/���El�.w�_�C�+��� r:�Mk* ����{9z7\~�{\>��R�@�\O��������M���	QOXC�j���XR2UUL�#'%?|�(2M:M�ş<c1Zc~�lI�b��b]�@��` �@�6�/
���*�xf9�1c�ĳw�x���:�����~�dxF��v��?��"*�-�GB�붸�)�B���X%>����!�?���ڭ#�[u\��|����hd�|&,�q�5�$���~#������é7"��j�{c�� #����_gs�Ig�^��M�-�h��8�͵3���E�}�tXvL���3�	w'��}ȎrQ�>K*2������I�}x�>/�׭�����4fe��V7��1<Q�qP�7}.�4T����5Q4��wn��y��if<�5����FDJN|�ル#����2�Vj��Yy)�ߛ\�Z��	��D��y��ɷ	�-!�L'|�[�X���oF�G�1��֑5ϡ��}��P?�b��3I��+�Ҟ���5q���&��]l����)[�6�uK�����ƌ�)T��/VR�2s�A��<б$�E����&'�|q)�W�g�|3#v��j�DS��QXk�]��=2+�I�9�_\���죵���"$�����R��
�$�ƽ6��w�sJ��0����Ou �?ω���Zȍv�>*NxD����ѧ�$R�,�L[B
Q̿08�.7!�Z���Y���z,s.h�y2���} ����2;�(�3Pi@L��F��ʈTeıCy�u��Ip%������kɝ�Ѳ��X�~�)���@�.��7���]_VA��5�����M��+h��i�D�ieR	�ŨZ��9��e��҂[}UG0���_��TE�����HW���NV;fd���;.m���<F�BZo�#\����L�7���Ά�-R�çJ/&�zVn�:�ȅ��t����t3�%�*���p!�=�zz(8��	�{���\�~|dyxK�a���v5�a�c$��7\����A�|��Ṵ������%H���X|<�9�=���S�S�\3�
���m�f����3�n�_ʶC93��kV��0(Q8��Ѐ}j��XS�څ�K������/O��w��p�;��|b�E�΋�:݇�ᒈ�km����Q/��7���i�	�%��d)8�{��er~MbDC���0U>6*�� '
ƻ��/̯C`��J��畎�8�wd_xN��M��0c��7YE�=�&���4i;��q�8D��Xݮ�,J
�r8��O�0y���!�����E��5���U����@���858G�7a�hmdcЃ~�(����lh89���SdKd���ڴoX:���ˊ+K[ټ@�.-6C��0��o�l��Dk6��V���O$^`ԛu����G��@�� c�
B>���j�:����Wk��X~I�x$�,���0�d�3�U�(��_3k?v	��^��x��<`�a���9�[��n���~%�.�*7M5[ɴ��%��y�+X��"��=G�uڅ��{�/�(D?�p�Ѯ.�/c�}�4;�,$Fasn�bN� ����Vr���1jI����]Z�Hư<&���y�dE �y	�;Q:K�0-`'f'&O0	W{P��ޥ,���ɞwc����DG����Ff淳r�Fޑ������Rl�����
I�' �2�o	����8�dj~�R���7��xw�8A:D�3g<j��/C7G~��\��:�G2/�gB]8���\L�| �+_�z�%�w E6���;������׍��"�je����������
^�7��9�� - p�l���Mŧ�:�.�i1%�;���;�d�d:�Q[()t�@�� �ϳ�5d��T��o|O�_HB�_`��֔-�"��������Ї�?�,�\W"��s�~>?O�y0�O�_Ⳮ�OZ�i~�ߙ]	%}�����3��7�jɋ}�zT�Ó���,}�ˌ�BGPm�r&3�Ӷ�T�=��Ơ�@�e�w
�>%�L�	hi2=����%"+���*�(��>�O�/��@���)og���⚥���NG%��R=�B~}�j7��S��sX�{��=��D��83��D��2�߻�"D�~q����ym����ϲ� ��SA�|�6��c�6낎���Z*�YE����m��6S��t��z��1�P��g~�y��
�G��<��L,ȼ:�.]lЁ:�_��3�uU��ʷ�~W�P^��C ���l�Ʈ_}�<"����H����ν�h�]b�H4O�ԧ˲�����K�JLF}h�ñ~�B}Ug<�b�HV�R-�sk�N;�b��Sq��=�L���m�oIR��^��T�T)��cP��-G��V�a#;�����Rv�k~;W��`N�w@�Oy�{	'��Q>(��-�M�ڴ�	�R�Y��AņbOh-����+���3�8N~�X';'�\<������;�a3g�����́��lA�z��1~�w�yO����#�-Gt��iSଽ$��xg	\�1+�L p{l.�D/ʯ����yԿe��~Y��X'�E'ر�>�����[�@��q6�T�/�^�f�|�24!�Tl"R U���������1s�C�e�<<�v_�ۅ�(���5?!�M����ʹ=˖�׽D�;'�4�nH���VƤ��k��^��r��O�/�����u�k#��T�w�L���
���fs-m!��Cm:c3��� ��i-�Á�i�T3E�X4���M'��m�]zw_�v�9A<�11ƟuS��w	��$��:8����F�u;&�#�Al�h��y�w��~�D��~Ae�����Ǌ,L��d׵��6��K��6��qi���.`�OaQ�U��j$�u���kQ`kR�8jW�+:�R���]Z���"/	����/1bS8g�}�-���+�4a���b� �!�+2�w�|�Q�i���G�꿧+��$�{D^#"ѓ?�]2��:�#����-�
�6�j8E����z9x�o=K�9�T�{���ͳ�	�%?���O�����*���|/l�2�>1���+�Hys}�\u�f����H����1ز`���&���S�."y�IM�iH�P���Ψ�D�˷��v��V5�RB/4��/�Z%�ɌnxLT���>D
�t�&����Qlt*�S���1�p�ֽwd�ڋ�p��r���zn�����i���=J@�L�_�^�0�c]�"FǙ��i7>ʡ��+��ǣ�7r�ݕ�k�m�\|��'�ܪ��ӗW��1�����<�ۤ��]:��\ #r�����b�rT��D�Kq[OL3M�V�-��@�\]� '��h����g��K�3�Fv:�y\הi9�6ۦƜ���t�,?h�k-]W9���0�=v�kC�y"C��a4��&@�~d:��PmT���\�pMu.�����3Y��Rrȸ*�j���j^�Q�=�F�ׁƟ|b\�DNS힋-R�׏>��C���`u�p �r@K��sC�P��sN|���?k���0��c�8N�L���
���ko��,NR�n������Gߖ��������^;���S�UI�'o]w%����g�GqLp@�%��ꚬ ��s#���(b���>�!��<����IQ��p:�h�'�apAN=T�����W�������'��m�B�wwwww_$xpwY\�-���>������7Us��N������w�y4� 87IY�}2O6	��(v)rI����>��϶�;�.|��0�966�w�`U�*G}Tp�v)�n �?Ch2��2�D+f�O�#�ԙ->��9_�?Al��1QE�6kQ],f�gi�����;헄�e;�Q���7�����5>[���Y�6��qno���|@��� ��<.\�b�#�6�����^��6���@��&������@��L��2�H�WIe��6$�p���E�e�F8�/����4��fM�����.�`dA���G�8���P�H�O!��P�%���Bnu�ξ7Ւp�ZpE�?��RI��ĳ��jn;�X8���-���@��}�����l�)��m������8
s_.$}Ȥ���(�r6�e��G��0_�}�M��Y`d�vR��f�f��f��Q��ŽT"���Ԕ����r���4�h�<���I�UXX�"L5
���e4�[�-�m�t��T�w�#ÊJ[��8z��f�Y0�*��1�E�����dt2� ����X9�7��1�t�0�x4ƃv���;�X�+N��HE~P{|�cZ�KN~�ts��c���,���A,�l�lh�D���vl>q�Ķ�����Z��"+��B�$��}�DG:t��f��<���F|���c�6��Ӌ%�&H2��G��w���`�b`����D�>�,|,��_�:��NQ9�i���*����!�Ͳ,�Sf
���b0i����*e�1�9��(.I�m�y���>�g"�s����5}�2��{�_�?��[~�*���tTq���~�'tH-��;sG���
��k�1���d�77ș7sl�uh�%�-�{��&f�!m1�e��ܖO\���չ��� ."���_Ʌ`LOC�P!�^M�0>����0���
s� �i6~r��Y��_��'���}0y����Lý�?���(ួ4�����n�x���zO~K�6b�O:��čo�<�[�������0)z io�������n ��?o��&��H"��_����o��)�E�KyG�O �����e��G��sU��V�$�HP�L�̜���.T^��U��oƦ@o�f���G(��W-�9zf�ɿ9c\7H ��N�+$���i����a�DT��@|i�`��ca9��CmsA�o�����c�w�L��B}��p£�`f�߉��RvpIs1Y} ���c irWø�x�(�hד�I���L�ޙ��[�e�t�ΘP�d�#��;��q�#>�+�qO��`�s��b?D	�%;�ҟ`�2�a]���gNk_p�5��һ� �ݐF��f-��?wP�y����9��S�ɱ2=�0�T{*NY�p���vA2�N�㟑��T��Eu[t�mӎSl��b8���`q�2�_e���̄����R$d� ���]��/D?>�uJQ6WH1-�lx�P#x�f>��'�ꃌC�@C(\8r%?�={�>��7�A�S-<P4Q�_�[���>�Ge���>R�
�yt�Ra�G]/�B�OH�.��=�`_1b��R�2����c�-�W�Ϳ}��Q��86�_j�?����-��W-B1�N����*����s��_��U�JaWR�A]�1 }$ɼUWt9v�>1{�v*s��
 U����.0VA��ӗMU8��qq:���?/����0O�����*�I,�n�\#��d���+������֒���{�}�DPA=�z�J�KˑG�H�]3�+&�t��e����'FS��U*�84ؕ�+�ڮs) s�M����:q��Y]��K2#��e�������,��c�_�K��N���L�sa�7J ֥��#��N��� ��� �n��Q�0S�n�#�KI���@�����ԸI;2����Ԑ�/5��ld���
11�~����E��p�}����.P���qL:��}#��$��N�������W�o����U�[����ng������1�2i�d��@>Z�R���R�p_q��JSd2���'�^Gѹ��<$`.����8r���'�B��A�N�:�C��S?�`c��f�mC��|�x����MݐG���Q�F��X?^��i�E��^�V/�6����b[W���F.n;�,6�����/�.��?D � ��^��4Dm�H� BZ9�C5>A��q77�;�ڑ�:�y�y.����Ӧ��z�=6��В$&�?��b����.@��l�h�$@K�+!����h����Z��`��z����%dw&��o����A��f��9�>4$�0���̐d�vsq����bc����U��jl�z��aD*k����L�toe���#i>l���Vx��t�^m۫ۚ�9�c,�d���GA�?���9���A���QK_`[�Z��q����+�1Vf/�w�9x��*?T�(�n� ��������<�W�]������n�QI�M��Ư���v0cJ��y���OJ=���^�K�F�D�ǔm���;�}�� ��V/�gK��l���gH�ֵ�<��A@�p�TC��7/�y~Ȟow#Q�xq���Y�4�#�����< �G2�p�Ġ_
����gc%.|��]�F���L�U�9{h~��L{4G��_��o���� Fq�����f�h��h�o}���_d�1{?ްmCF�v�I+ �]�� �!,<� �.����dvZ�w@��m�"��t�dW��W��*�Cݹۯ�ݭ�>%�E "bM��w��BTP�wY.P=5n�)2�T�����b�5�m?�x���w������\���;������-B�����\o�\��  �?[E����Ϗ���nU�����I�I�p��ئ�^-��
h�jH�4���GI��<��%{�6�\�)� f��!��B�?�2v�S���0j*�|>%�U�����;�ݢ�{�*LDL���n�HK�搠=�wĶ`q��#�����C#�Ҹ���������i3{�5�qED�����|W#��Y�#�L���q��{�1��+�=�y�֟�cJI�=X��)�r�`dֿQ�)�d��=�3�%vuc�v����j�"��t�s�9�ɚ��q�/}�2R�)U�VkD��Nw�+{ ����4�>W(}ė��9��5��dQ�m��5�U�Z�<oq�cc��B]א��p�M��j��DPNoW��J���{4�@�ej���Q����_F/�U�J���M����&��ؐfzj���	�(*�&A�;*J}��E��ƛ�f��̅��~>G�����&��|�:����g'���Ȣl'x�}3�����;.x:d;�g�*�:���|�y�p����sZR���Ѵ�ar)�v�
Z蚌Y�9�R��=��8W��ިu�3Z�p��eÝt|�\��A����`�Uu�X��w��G���/p}Xl����_�]����DU*�{\�3�Aq�]Ŕ�/eX�-(�*!�;t#V���幚�S�pM-_;L|&��:{r���<��"�Z�G!�L#�`�h���U����
���n9�� �IGl(�f�PGnq��UN�z�h{��0h��8�D�+3�{12Gӈ�ʠ��D�Fek�P�c�����Tm�əv�^T	�f�>��v�C��,v~G'�,�ڊ#}�Ө����5�IU}$�(_$�TF����/j�t	�	�r��<�
��j}��;�X�d�,יK��⥀~�G$�_���l
[�5=9N�٢���t�D~�/ӕV�� �F����ݔ8Ov6q�4Bi�(ЏG*�3ؓ��־�4��d�m��V�U^�c]R�^s�Q<+|�7��M� ��'�|�m�;3_\�f�g���s��0v�c	�fsy!��?WR��.6�8����c^�u\��=I�X�-�4���pN�J6�,���}��֓�1sk~��*����dG���Z��Y���ɏ�+(r�X��r&��>�߈���%#h-�}$�VQ{�8�C�� ��+�!����b�Ǿ�U��f�8G�Hr�4��6���J�P�p����o/,���a'�h�\�R`v[ELXb��ev���	��W�O�KK�Nyp�i�e)�.f/`rE=�y�[�<�i��qiO��&y)Y���/��jL2�ٙ�5�^�9�[)co�~+�֜��*���oq��F�J ��ؑ��*�2|�mL]7��&�&�+�BIZ�b�8澣�M��B���F/Yc�7���d!�%��%��0g�Gd�8�9L˗¹�I��}�19�Y����s	K�^X.7Q9�0�1�;�"m�������P6���[��Jb���i��麏�z'�"ȿy'�J�N�����i�XQ������MH��<57�w����_QP���X���sd :�{���ݧ�L�h�5�|�jD�p&�(p��-�	Ot�%�@)��5
Z�pΥ�U�p��(���s]!�E�N�s���]��v1.ؿ]�~RBk�Fߖ�є�n �y�6ư(���"�/�qKC=/R�^gW]C��7+�v��mV~���!B|��.c�)���������.�U���.�,�ok��r!�����2��z�ե6b����n��Vj�bl���EdJ�}��( �`���}#�KW{]ֺ%3�چ8�K��1���$�4?��M���Xv�f��K�m����8�q\�XJ+��͹̦z��h�`T�%'��c4��׵e�I����'h��S���ѯ�Wr Q6��m����R7��ϸ�6���y?���.����N��,�6n#ptG����5m�<����a�_��Qn��rF��,湌�6��9;�,c>q���B6j�8�?Q��� ����x��g~�_F���r�B�  ����A��F�+M��yeB�O��`.1F6��S� V!-i_&�*���A�f�)݊���ݞG�����F�S��;%-{!8-�a�8�餮������P�\���P&����n~��I��j�/�`�%�H]2�咂�.�<'�0��#�tI�T���|���H'��[�X&�i�8W�M���~3��$�Ex
i'jk �"��s��)k߹v�^{9��!����P��Ln����R5����MayX��1lB��K<sI'h�J�<'^�s�=+�'��$�$�y���۱�'f�I�nM�J6�J
o�l�U'�L���k�HZ��R��&�"���}����r�z�>����n�ɡ�S���0lp���I��9T��L01�i�í]�E�S���s��s�i*ʬ_>�[������Y$��"u��3�#�.���}#	W��X��⇒6��9�(G�v?�����K���V��P�u��+\Oo4�z)�>��t�!��_�q�ID��̕1��á�#q&s:W�G��_�	9�]���R��| �3q��:��ZNy�f�a�S��A�T�ݔF}���]g��L~]�	��PT<}���	oh4��X���xn�v��8��n�,�hoɵ��|�ZXDb ���Hy�~�s̳��ƃ>�3�@M�0^�0]f�^��(��y[�ݒM��w1�mvA8.Rn���D��$$�w�o���mT%±�h$P���G�e�A���#ӝ����h�?�QXB�P@�+�{!Dx��F�Ͽ�)]�'��He�~8����VP�%�j�h��z�ʹ�E�2��e�+͆lz�mLa1�{M�Ej9.i���}���0wͥ���	#d���Kj�{t(�͵'X�ߒ�i���a���b�&%TB����w�[F�Z��T�D�Rө�t��?dl�W�.ee��pkT�p��}�-�����}ɩ	�M��.��-{g��3�����T���+�r������qѾ�g�זQy^|6�e�I���Qo�0`��̃te�0H&�v,X/�]g01l�Y0-e^�%@��\�8He�+G�Ҙt����)hO�B߶�n�&� ���2֮�s_�+�U܁8��ʹ1�#ċ��� ��wtχ�D��[@��r����Mw����|�E���?7�8Fl�ў����=��n���c�6�/��d��*]�⏩��8��=P[�-���&�Ǵ��.�0�F��A=����YR�q��+g݂�i:���*����Ƙd�}cMTp&Rl	Z��Z���b�px-�>U)�`�)T�zf���� � ��4�j�%WKu=9��?(2Ky�]�I�'r�>� ��l�xJ�K����� Ͽ�b���.�>�mq�g�W�=�3�e|�����ư�;r�B�3E�� �9k���
����)@L�sTW�������	�4ݍ7���G%I��!�{���!�$9�Wuu�󞌟?)#��Jئ�ttHN�7��-ҽ��1�����m���y#5�7>+�gZܾF<^�L��\���5z��
�w��p6���r?=T�N� Ĳ�~V�h����:�&>����"�0�v4@|C�����L�rX��o D^����M�y��flsz#f�)�뿄i��a�[b�%�����|���B�i�䥑OB#~(����b�r�w^��/���{���9E�M�{�6����s��쐌�p����t��"5�F���h}�ͥ�6ʅ%���M.˟��{��W��֣���f�y��k�;���[-���v�ᦱ�H���2���pA���{�>S��}ށڍw���x��^��9��!��ƀ���2����yD��eJyHJgX�,i�R�	�F��O�j�Cm>�C<kc�4��������a�'�-ԡ����Z�y?�5A��J�8��u8��|#���A"Öo)��ح	���a ��� ��Π��<�%�nڪl 6��l��3Cs��'�g�)+F��F�|�L�������&��$wAX+����d>�V�P�<%�ʎ�T!:���]"��w ~ZC]��K��=ДU(齲�~��,`6JO6�Mj��c������/�Z��iz�<����o����@�G���$�lGt��5Q0[��V�b��̳Jݯ���N�Qb͒+�);;�d'`�|�-Qptz��\�"��è�x���N\)f�0�2�7��H������/.��%ל����^l�_q�+1���3�ڴ�ǆ1�S��["K���缞R-m���p5�]���>w9,BEt�PF��/?"F�������V�/^��e	z���L�r���J�)A|�(��t��	���N0Ԣ��t�L�f�9q��L�'�s6�<����v#��f�	;����
��-=Pg#����R\mɈ&׉�"����B����w�%�y��	���r6�W61��9�>x;b:��h�[��C�$�@�A+�{/qZj�l�� 
�}e�m�\����x��g]^e~��FYĮ1��B8p0�I�<��u�����ߋ�����/RQ@�ڱKU�}�~��X��/~Fi� t�;�>ڈ���oK�Jcp%�;��s7�&����S��զ ����
��Ј�#�'O:��֩��+gH۟���S�Lt2��	hF.�
� ����G�5}c��1�������Pv@��d(G;��]�$q��F�D���=�ձ�t����l"Z�o訌�\g(�'V3�*�8���(�����,�L<�4Io�!�S�!�Ǝ�-���^l-�,9,m��1�L��i�޹�g�G��[���~�=�oR�]e�85_���C��)��;t���3�YOf�ڍ��u�~T�흔�R�x�XjԖ*��p��8ᥗ���=�F�1"<�>�"/�9�]�:�Zr��w������34����Q�����O]>��!�視db�"�ti�_��[d�[/�i��rYeo�yͽ�<�}��󏊙]�qx�� ��hV���˧��Y��a4����9�0���Pi�(�}���fL���m�R9�X�QFʂ�xE��z����T��H�A�-�̖��ᰡ�KȊ�e�\��$�*��;g��O�R}�:�X�v�-wzK��q'�|�H�=��8.K0����ؙF)9�j�ː^�I􈖲�m�ڵ��*ֲվ/-_W)�v8V�W+�
�+X��t~�t��$%Uy�ȹ���&|�����d�A�)�(M��b��?N�o�?�յ���-�0��<�\W��lr�@��)�{����v�FCZr��}�4��b�����*�˥��ϒ�;�S����
�!���p����)�����! 4�{5�kD��olkM�� D�K��]�rD|Lq!�ONC�HrQ�ge�H�����j�T��S ���Y�ͼ�zه�°���y�(��}@��.�I˞���#��+��?'{U���"ObC��DY�/;���e��������4r��9����D����/��0�j�V&��`��)b��,w �)d��4���`���[�o��D���>B�.k�o�j�f��l���9�m���������Dhk_�,&?%ە��`kr#�z�w�ݓ�:��)�kL ���r#~C
���R�6
i���O�=����9����B����'����^*)&k���9���{���E)�"aAY�xA\�k�I�g���e��3��(�t3&�ۿy��*��OCi�N����Ȱ�.;�K~gX
�O6"'A_�9�}:C����>�e���\�G�A0"�)w^G����i��D�E�|�M���Vk�v�`��׳w"?���B�_ō1z�-�r�#6b?5���R�=�gH�0^kP_�9�"���.*7]ơY���<�vp�r�i)���ѻ�^��]ى3���-¼����L�O�:���4T$'�^�����j�9�?�J����]��T�a��zC�f���� �@ޭ m8��L��O{�<|�
�Q��d��.L���{��y��r������QF��۠{z:<}�>q�/�g���RH��	*�v��]|溉�m�;�#�*���FAA�z������ ۉ���-���O�e����t,29vZ��r��OC������G$�n?��a(&��ulɟ��w�5��4�٦Iȡ+�������\�
���<���
�Y<��hn��2n��H��kt�/0t�C:���T�f����T#�O;7L���3��$l��l�x�J%z�yʵ9CE�Nos�0�~IruJO�fݍ\�5AC��2X�z��AhC)��Z�^$���<�?�^���N�P�O�OnzO7��_�<jA���8�zi���!?�^��p�,|�J�*cQ�l�I��ɖ;z���ʰ��KA0A�a�O��F1�q_��tꇚy���#Y�Dbc�v�[����s�Ac����L�18������4.V�ȶ@�	���.0G��������n˒B���=;��8S��E��ZT"-hv���م�=�%?G2�K;���"�,�N&�#9��_�)��c��`-��;��| T�Q'q�{��x*=䧬�V�����A�X=� �B�9���	��/�'�f�=������?�Y�>O�t��̮�0+��D�?��a�z�n�f#o��~�#��P}�bSˣ�`ã�P����܅W	�{�&T�
��\ϳ$��m�E�)L߀ǁѨ�8���?���r�qg��ec�"��J�/Z���~���^:�Ob
�2�zv�2�� ��ѧ`����T��l�iޜ�����&�i}�*���Od�&�����
�0e�D�g����{��w��#u �?rJ�K}�GRy�ض���;ͧν�>�?�����J�"�ꂋ�P� ��� ~K�*�x���a��4p��w��an4�6�ӎ��?�A�%z��޼Ӫn-��o�"w�OШDQ2�UE��<LL���ѣ�l�'���xO!�ù$�֋�����aCe*�
0�a�Y������~><͊�SY�����C���/e���`Y��^���j�� ���c@�����%.�:e��}:*���R[�P2b/���P�X�>	��d���L��(�ޛ�u��q�b�9CA���5��q��`fOuG0�0�;�{9�W��N�R��̆�Q/^�n&N��~V@&������-��o28��A���x�D�p6m�_ϫPP_��9_�C���b�bҿ�����%�Y%��$r'�r��T���̽�f@3��6�E�&׬*���&�|��7�|��6���L8L�N���1���[�-h {kneZ&^DER��a�/R�rH嫚��b�!���R:�ɢp��Il�K^Q��m,"�zp�N���\���F��Af�U���V�60��M}$��\F=5ګ���ʋ>ߩn���RIn�N0�骙:Ür���~�g�����"�.�C��=H"G�O:�z7�Cr�H�-�XbjѦ�����HE��z.KU�1	��Qڭ�����O/���'q,�7�qv~��ky�c+x�]+��?������)9�_;שn�M���O�)�J@[�S�2���:�8g� ���L�"o��6�Ӌ���EM��U݅���s�&o��O�:qqS���z�\QL��MTҙ���q�S��\��jB��j��Iu���5��\� G��^�c0zF-��M�IF�GTJ{����B�[%O>�g��vD�Ϥ���4�Ba�2yl��u��HH���50s��V)f��*"�9�������,�_�
&��IQ7�֐��%wz����<Ż.L�W�3NOR�t~�:�H"�t��x��Ts��ӣ|���4������qۂ���uQ�9̬#�尠<p�OW����6�$��u�>��jOG�<�[�|4ߪ��E��t��8K��)��R	��`y�uV�B�V�k��������"�0��������En?ه���R�6	6�5M�4��S���j��$R�$C���^��O����b�qMK-�ў��M�x=�\�l!H��d�g�s�I�`�]���<�_����}����O3#o��%<^Nn�0��"7�5�8	�|�x\ܾuǇZ�if~��a2�J� ���e+
��+J�ś3OH^���ÿ#��A�\�m<���f��®���U����J�.g8�%p2����|-����B9�����fA�ٔӯ���B���I!��7��I�z���P�}�����]�vǟ¼��vc\܀��N6�&���SB�_��ߌ��Db ��08�� ��L�1t��͌$���q�>�$��|��;F.#��Q��q��ÈT��$!�eس]�}�͋=���*�~~�����L��=%�\��w���$��
������q����:�X����y�,��,ob����$����+�����jW@�I*Źc �Jׂh̾�� 6��h�i]*��T e��Jq�~�&4De�J�m�9$^��|a;�Bn��36�Ν)?嶢8��{n�;˟i�sA�^�L�����g�!y��"v,0�~���>/��q\\}d2|��$s�i����fp4XY"�����=
ޞ�c��6�H�&|#\�9���Gj�O��͕:�~?���]���H��{��3H���.�?���Jޔ�B�K1bH�]ݖ��$����?8�?�>��f�:mX��6ED��
�T�pܓ�N��e�5��WW=8;%r��� ql~5���L�0��W��u���oi��u��Ao�ɽ����v�1��D+h��S� ��<X��rZYG�Z�˨�O�V��I�n�F2��We���!r�t$P\��V��\u�m*0�vT�3@�q���N;-\)F�A��o��6/��v��g����Y��d��yʞK�˅��6A�����8��+�F���ۆ�'|���T1G��P�X������֎��8����O1
�iǽ4~�AJ�F�3/W�¸�"�:*Q듋�'N7"��ۇ�e+�BD�?�%I�͎�m�/e�{k�VL��ʋ���q�i1t�oeW��g��E��z���v�z�װ�,)%gq��oGn\��7<W��P�Q�Бb���R���dٞw����S�\�&�Y�w1mv�5��
�7�;�#td&H������G ��\?������F+����A1bjj!2>����-'��g��N8��]����l�5����m���[rJ>�bv�ލ��t=(�o�6��rOKc�Y_#�^�J�&3��>���ʒPŢ[Ӈ��p��C�sU��X��)��JF;8�I?�݇���6:>����U�_�g����\�=t������9�B�_�M��[R��e�o��I�&��/&�=p�÷�?~��m�̊��<y7�[�:8x�!&_��]a�U?;�e�V�ޜ��jA��4�O1���k�C��1c�=P��#����x�5[y4����2��ƙ�N�d�N�V����ͷ��՞����ui����[m�W�gaj�AFϧ�VcA��cf'i: P��&Yǐz�tH�9eLd�	{��Iu��em�#�K6Q�[_�iR�E45�P�0l���.V(j�A��/q휧I�R�w"7�;�ߞl�M(��d��&�*��GpGAf;� [� P�m�MB��Og"gU�Z�[����a��za��E&S%�7�O�����ӱ�Ф���N�L9%1�l}�����IЮ?��]sT�Ә�[6��u*�C��e:������G�=�
���ҿ|�%\�P&�K�}2�9��>�����O\�:i�Q3<p��{�t]HD�Qº�t		��X�� ��[oV�ƴ7�T��k�J<�b����f'���v=�x���l�ǫ��_Kž��︸_ܳE5L,
*խ�N�x��ͽK��@���)ȧ:������'N�����r"c�K����sԥ(����[�'�Ӝ����U/	�AJb���C��T.]Y�K�.I��d�oη�M;>��w�>���Y�#���0�������vu�<7> �]���p2��}5��<����W@���7k,ww�DH;��+�3eX�[�T��]��-�!�����쭀���~�2:�s�3�s���� �7��>�t���^��s`��c=���<y�2�&�U�����0Q�_��)\�?y����a��	W t��b�oӡ�^4������%�~W��G�o���pʥ��,����;1�&�Jk]�|V㛭v�VY+U�(���oa�����?��Z�hp�\�g��BJ�p�Z�P4��C.=��jld0`<ӣ��Ӌ��rĜت�9r�5�ȴ�P�P`sV�]���Ϟ�:����>'��
q�&�aZ�����u���l�&ߣ�p�@���ʃ��%��0$$��$���|�����l���܇KZ�(�Vj0���h��nFf�(I���T�eo��s�*�1Ѫ`��P��kta�n���39�Lz��bJ}.]��8��6���ڛ����t
�K�g3�N#�� W�M�9!�/�*�r��'���idc�qr;�wݏ{�R�����\EDĥ�]�z@H�~\���n��UC���lK�Pطq���B���L!,��H�6�y�&�銡Fn��V�P3���5����N��%=vg"!�d~ap�^����>
�u�|w:p�c�-2�,�tg2�w�)D�J�ߍ� ;<�Ee�i���ΎM��}��v����v�-}$�K~�7ޟ)��Қ�U}����Gs�%������Y>�,���1�;/���.9I1��~�������z�������;�}A�cG;!��f��7� Y����n�论��l<�zvF��ji+y��39��g֙b�	��D�+ދ�i�1a;�-��B� ������i�U�H�G�z�O�c��m�m!�w=r�Т;�Kƒ�����b~�I��Jp����K�j�o[��^��Ͽ$�m_��l^��S��j���ٻ�L�;��FF�U�ӨǈA5�q+��Ie:%�w���_� ���+��F|�p�f�-C�E��"���X1r����	(�j�mw-��H��~�[H����6�/�6�3$t�x͊"��]�^[_���5%�����s�G�S���>�j����\����;��aRޝs�Z�SL$�$��Xl������j��R3�u"���͸S��Z��22c��=�$+9�7�;�ǁ��p��]89�K]�#�7Qh/����L4�ly#����[��"΅�݄�|ڲ{~����~u(5VCT��b�vי���Lsݗ�ik�������3��R&���W��ؾ;XԳ�OjO4r���v�r�6}�WO��xA�'d83گ~�S�q6q�R�.�5�]���L0��f��o��<�!
�:VC�4v�����\e����)<�ơ;����
� ���ec����]]�m�j��>[um���p�����9�v6{	f<�fK %��=}��{7��V=L&��ƧOdݎ�t��<;�g���Z��q�>C~5��k�'a�~f�f��=L�0��A2���9Ͱ�z0�F�d�b�4Մ�(�ɶ%L��bi�����]ϯ�GRvpɠ^c��z��@ظ��᱉�39A�Q��Ν�(����%8�TqX�PZ�&U������&KO}dZM�/>A�E�o�o��;�O�h�*������>�!��5�}�V0Qq&Ŀ��`j��6h�Vl����|rh�?!�R�=I�p����300������J)1X'�:�'BG='�� m#q^hG��<v��G��(�#�������8l"NUͅ���<-|{��m8����ΞtL���8��(�+wV�>;��՘M*'�lb��ӡ�j1�a���:q���]37㤝f�ե԰�g���|mg�����h����A����o�n�C��V�,��JOö�GPS�:��$�DU��J1�B�D��E�'J��
��`���ym�u�}m���C&���M��m]yk -�e�z�>[�"+r��g��0#GO���y��e�h�g�AԲ�Il��b��X�:���0��+�����yf��+-�-�GX��B�C��L�B'��}eU@<Ȃ�r�]����,�ʂ��2��V�y�>b��N>�G�uw83���N~�/P������gu����(����'�+JJ��wr���L�?������&��F�9�+�x&~�b�f9����JP&�6��#KN)s�����n���[;�hј��ݟJ��~�C�T;���m��c�ʟ�R�g�5#si�'�;2�?я�N��&#�lՃ�n��>n(}�;=�+E������C/��ž�]B��ς����1��xz��α�_*R�拌�_�`s�*9�5~��?X��ĵr�I��;a4�A?ns����0驹R�`�Ž\��͂b����y�������X�F�uDS�mX\�~�(�G;�͑��B]Bv��"�`����%�EVQ���G����׎{�>��sh�!�;�Lae�ߧ�R�I��9>�����u1돮a8%?��^��oTh�Y��)��K(���㴪c�׸�k4���*!^�G�	[��7bc�@�?J��{~�~�.C�P?�В#X��7
�q*�T����%�Y��v�'�`�������Z?��s�s��)Ėa>��S�j/��`H%���4D�j���1���u��q��b��%��z��(�%���t�,��P��ݑb/)�h���:�Q5�9��lH$6+�G���<����t#�j<��ǥA?�^�&��j
�	˫��,O?п��{����&�ވ&�3{}o��磗����*`@,p�Y�CjC�Ĵ��!������Dq�h��T*��Lٮ����P[N���Q�j�! }����|4�lV|�� wh�ϱ�7>�	�ᓷ��$!ŏ�$V�R�Y�7�����x���b�(ۢ�u�n�+68��:�b>ŌR�U���S����xoŠ/�ZH���7P�e�ۇ)�T[)��s�MB�������G9�(K�E� ��:�H�n�����܅м?<ɷ�Η¿z��F���k�6�+b;��s��I�E������
�L}�8��G�xZ8ZfI��b�������#�����Puq��#l��ٽ�<��n���C���_Bޝ����(}>Z$^���i|��sW���F�'��q~�� )՚l���dD�P&�Y�oZO��a΄J?W�`�`�Xw����X8��D�5x��9��\�h΅��@N��WtWέ8�Q�#�Z��\lw��!o���VvP�>㧰|ɾ����;? ���FMO�-f3���Ar�q/�lX�\��ժ����ڽ�b� e���ɔ�
�x�"��u�JH��} ��Lܹ���DU��;O�q�*�$�ּݻ{������nk���F	 �z���"E@:�)R!қ)AzWD�)J��I��PC���{��ُ�>�\s���bf�9���=�$6{��ɫZgV�[��.�8���8��X�>~�Ux�7��DY��?��-�8� �bZ�)�!_We�ugK��ܩ}��=�O1�7�q��a��*��ЏY�xmo�%}ys`"��I5��^��^H6/�u"n#\-$�l�n�|(k������;�/�ǻ��u6�f<��V�~v/p��z�'돪d.S�v�h��TE�U��jR���L���O\Y�#�M���	`��d%�r�wͲ���y�+�v�D}�B��Г3�����Ӊ��Y���8�Kz��e)n�vS�2���M�]�9���.�0���+eF\�ɛ�������Jz��]�a�׊��v�����~�My���NLݏ
����U2tS�~�&��,��1�<�&}�~I'��Ȁ�����f�P���K�fC�(��O[�0� �	or��c�8���`[�k����!�!Ռ�>�x��<]4��џ��G3o��h�f/7Io� ��?�ʸ9:O�(����l5���r�7O("% �������-�~��">���wz��c���m4�N�|�s����6jC����`�����;�'�\{��o:����z�>��Ǌ���X\���W�4�z�c��B����̿yb�S���1e��-�*�)c:I:/��m�����za[�, �7*�2���0�'������4��д_�;hGWi��k��()�I;�޳�y�!=�5̶i���Qj�}�/���E?�8�c3�~y�m��]� !��g��v<���y��� ��.��g��9�<b��]m)l͞�2%� ()���Jbz�+�+ί�G���9I�0f�������o
���������4��a�u켫�sO�������&7F����^�����x�閎��/_C~��)���l@�q�>f�k���"�#�N��r�m�J�I��@7_Ȩ*�cj��\�/��KZ[�m3s�e�����v�Ikh���l���a?���o�t1�Q���s=R�C�O� (��m�X+k�a�/��}�9(���2W�_�)~�6�޹�����u���&�("�f����?��yno����bS�������r�?n]��TLx��CW/�S^$�G��^��G7M�W��g�Ob��~�'Au<���5��0�2��c�֜����Qո$�hG>a��+���ӻ��_C���P\tg\������;\Jfj��F�Q����4�#H�[S�z����@P�Hɺ�W��:A}��I��w�������
�h�$f.;���87��z&o�aS�����n)�at�t��v�kP��4G*#�g�<ษ��Q�f?g�>/8�k��u�_n�f"~� �:t�r���^��- �W1�f���ݍ���_`~<���Pib������8T-�:+#�v��S	j��"�/��v�w���
�����a�\���I{��H���Tg��_���lGjX�컪X�Ŧ-l[�u�0�V<���԰���Q�T9���B���~�����2v�*n�J��m��p������F�䬷��u��9Rd������gU�,~��s7��r<j���a1����08�$�qU9�1�=�?b�Y��R=}yҹ�0g���ر���:!w2����_���0�	��mNC:�������k��9{?��+���6�}��r@;�L��y���(�\N���W���'N=�����q>�r�S�z�Ax��x^�����9�ݝr�7��.v��wL>��͢��~�ym�zB`=Qb`�6���6C��i��#�O���3�ҘQT��Կ��YC�F (��k���y� i1����ҋ����b��L��;RB�!�6&�Y��@,�P�����ؖ� /X�^b��{�loO�6ֻO]�Ԗ�( �e����a�����iMY����v楻���ڙ����q��-�OP�����v���j���[��S�	��IF����W��b�!�̦&L.�i���L���iI#.|ݱ���F^��r��ڟ�3Y�|Vn�9G���R�a`��1��9�FYی(+���_<=O{��)+�a�SSI�S(��5e�����Q��F�d�ZG���`��g�ܪ��g1-�E��P�5@q@�~#3�0��W�@�] !���Xow�:a9!ee��1q1oζpһ,^U_���p��C/|\*��ح��-v�� N�����I���D�Xg�W��S,�[�d�T��� ���d��41zf�������H��`����Q(�<V�x`t��{nP(�����ſƜ����Q۲��ՙ��kE,�7)СT"�t/L�< ���]�����c����0)��:=Cl3oy�{�}	J��\�ªH�vT�N�Q����M�G��}���5N޼��`��G����U `Ņ@i�=�a�i%C�Cz�)B�99;+�w9c�_��������&LϢH��(�~�����Mڰ��D�'@����?7]��T:#��iH�Jt�B��/�1xWb�Ȁ�"j q_E�G��߬4=Ȑ	u1�tb����`�y�-��g=�O>g��m�!g��y� ��P�Q����0����j�������p�*�u���yR���g��=����U(&�����߱����[�r��܃k�d���Ѡ�g���(VU�슋0.��!G;��)]���e����x�	6�>ӓV��\cRe�_k8k&�9|�D}ys[��Z��=��G'_�M�Δ~ⵙ�*=�9p���y�ݓ�}�F��e� ��K���a���^$�v~�)��	�w!l�����|ζf�U�6� |����_3}u�qs�UsT��|ېE�<�x2I�@���/ݩ�F����K��W5�����gD����ӟ��^�57�Ͽ��=V�b#fk@��U��1�oέ�e�։�CțnC3�B�4f`���S�lC�[��w��1U�f���.f���N�0�!U|����1�Κ,_��iH������ͬ�W�yZ�~�.��a�<��lD��gŏ����_ԝ�Z]j�c��O��W����|���ӓB�M��]k)a���S����,��l���U�|�� \�!��k��<;�z�e.�� ���U�ē�Jz,�x�)������3������$S	��>r���©6�=�~j�[��8�o���B�ЧPg3H��v�a����̌x�^Ƙ�n�G<�?Y��!»ڦ��>cC�^](�e}�6dA)�%�}n�w�ak2N��lرTl���+���4��$A�<�ch K$����]<�2�̤FR�q��Ug���D�ș�֛��`q�  ��4�;X�К�ϛh>�D�3�c-t��"G��Ο.��L����� ��*�4���U4�䷭��X�/#���]�O8E�(`��K������01ٌA E���4��X�qJjQT��xR�MW��1�\څPpc;��ʭJ=�f��6�QQ���KO �r�H ���{�K�Ԁ� f��f~}ٗ�yA\BC�w�iO7rZ��@`?TSˉ���o$�~���J�$�N��RA�,��b��y�jit���y_���L�Ӣ���UF�B�&ӛu_+ ��ܽ!�Bc��C���X9k��6e��~o�{�{y�I�$�����D9��Ŗ;b��h{�2�-�����L��t����F*���r�����ނ)n�"��D��:�/Zey����a���F
��C��ӎ���W:ǟ�x.�o6�����.u�̕���������`��SԸ�f�1{Q{w�i�n�vp���.}�R�F9@�7p2��{�E��_C�Yr Q��w��)>ͤ�O���C�c�:>�:z)2�}�_��X�x�@���?��?���(M�b�%��)`{��.�+�������Z��$9�5�mX�( a�X�m��gaY�@"�=@`"��	'iR�{_��㶐�	h��d{�g�|����#�P��J�1��V8Ʒw��(���<J[r�]�ة�'�T5De��ѓa<�[�εJ�K���2hō x��G�Yה��ǻ��}�M�>�<$�Zl��=j��������9ũp����~Z)'6��F�3a̪Q/3��^4"X(�&~=u޽��zN���v��6��W�j��6�bȖ
�KS��1�&H�-��L7��|�����_MQ?8��`�f`��}�/`.H#��Bݹ9x*�;��i������@�[�0A����H��$�ҳi�T��6'�W<ř�z+���v��V+�L�0�B�{�����M��o�����CmNc�USC�G��$(��	�!��Si�
�3��Za��ZhT���(��G�e��x�;Z7�̿��VA��P"o'Y�q[o�j/����o��e�O�Q�U2��) N��[PE����Ům�U&Ʀ5��,$�t��o����E6S��_�w����|ַu�ن���g�h���3=��K�&�g��V���{���X�7ʱd��<��ʜ�	��qr
6�"�8H�q�����2���]Pӳ� `u�X�E��u�YaaRy��,ޤ��e�]N��&�"y-8Xx<�|���NP+j�_�H8B6�'c��'(|Xr	���W� ��:u���{~��r��;r���m�01~��j� $����v�/Zfդ탖�P�g[��"�Z�-}
TFTe�Y��Qϋ:;�{��0���_�!db����6Nm�]?D#:G���;_75����7'��<�L�6�͔>
��r�C��O�Jy)ѻ㦘�Ñ�0�F� D$	Ex#�$I��C�)���k`Gإ�\�g��<�-�P�8�u~�_�:#"$tyI�q��f��wh�F��'�&t3q��g"1�I�H��i=�������^��Y~����֠i�T]Y�� 0����=b��o���!.\�~ ��e�/TH�*�q8�����*���N��Z���Od>$�8��20q �gu���
����T�K�HJzV�*���>k�M`�� ia,q=�6�g�u���~9qtI�����eTE%����W��\�}<7L��%�����O*��W+J��h�O��ʠ�ݺ5m��7��蟯 �2��fB�,.ʔ����ߞ�%Z��'�-ھ&,-�ƅ���yL
�Z��ż>"2w^�t��UnH��p�>{�9�䅜���_�VV�=�4�S�+8�) �ܪ�XOeB�C�^�U����3o>�u�myKk۸��Q�U1��b�]�t�H�C��e��Ps���m���qǇ�|�3P10Y���m\68��%:I*���zS.W��C�1�Ү���	zx��h�?�;��-G7J�}�)V���:�Ix�d�:�S������,��˫��{� ZdE-ʙc��~�2���Ov�h�^��
���>��SX�B���S�
VQ��C�x8�g;ٜH�<�C�x�?�\x*�����C-�ۈk���/�X2��'x���I����k�"�L)�3(��#!E0-�D�d_��G���LI=��E9�����Խ�%�#j)��'aBB
�q��%E��b�o�_`<$Ib(B/��>�-Cn�6�'*�����%Kݎ@n�c�#�g�N��
	>p(��w�C^i�e������ў��s��,&w�}wW�൞����x����&�דаvt%�B.H� ��*ln7�=w�|�E6��/��jb[��*n��q�~���Ƞ�E&Z�IC���9\M}�O<w��.�?�W.��A�����=-$`��Nagp~4�Ss�'u('5U���o�"��ǒ~aH�	�
A�[��t�v��3��X���~w|�<�.�U��U���R�e�I4��sDq,��!��^���GS�͗V�)|��,*�P�}���b"�ɇ-�Z�pB���R[�t6�� ���ɢ>�k�V^�z��������c��'�������
��B���gk��r��Bܭ2��g�����G�*�}���^uI�Yn��J�׳����w;z\(�!�ޅcūX���$د5Ce5�I
�T��1��^,�7a3��7p^~���Ew|��%|�����
�O�׃oG�{�)Ql[��*��-^S�>CÈ�o��~�q�l�ɼ���S�,�>�U4��k�l.P�WЭ��DZ���ۉ�̼��{����t3OZ��;Ƥ;�ׅ��6z�8j<��	Bo9�s�*����l ,q�;�x�\hfe�u��#�|`S�1��:��uj�����Y
����	g��E�o��k>�c�}�Q��8MI|�hsLc �;w� �	�	K偳�~�B0��5�C�^�|�9���*�6f����.��ڰ�C�Wъ��Ӓҟw�Ӑ�4�RS����1�\��C���Z��{��ۑ��	�U�i��P�ߴ���İ���~��t���0ۻ�z�T��d�h��Ӏ��_h!v��R�ժ�pqn�&���GxE��l!�Rc�	��YZ�*Q�L�D`h6S�P{K����W��7뵪ĳwl=�!vA`J��-Hf�++�� �MR���\�+�]���G�� �&�����G�k�a=|����F��I�P�p�Ef��da�)ƹˬ��zX�6VT��|d.��G�m:�إ��AM揁} 0}�����Tp�}���,D��m���ԋ��)5Ng������k}��aۘ�Ɯ3ģRL���<n�����btV����t<y�ߌw&�&�����G���������`��9�:��d��#�@�ϫ
���Q2!ޫ��#hxm�~��;>zB����J�2��T<��!�,J��Tk�X���nw;Mi#D�{VT�j�M��E�����Z�Y����{:��J�f���;`0�����q��� eV�޷�G]4�D�C4"z��>3��!3�߃����Y�Q��� >��J���ҥ��[616��������W���[k!�b�$_aߠa��s��,�'>�}҂��g�����o�u!�S����I{���<��D�S5��٬c�4��R���:�@i���������:7���� ��(t��@�W_3�B�(F�>�^Ry��j�Ջ�0��J`Xdk�j����*�nR�"B�����q�Qp�D�P���:�'��a�z@H|���䕐ETd�Y]Ǉr�Oy10�m�ާ�,d�����R�7�h Rj�R[!���h�n�*^%��J�J׵��m��)��ㇼ�N���~���YY%�$�lˮ�O���_)f�*���6��������ڝ�ۀf���=j��նRmW��_�R͢2RW��w�?+�x�ΤiJ�6;��_�Z<̑'�U�Z��氳���:��Ӽa�3���4�a��<������Z�֥��c�W��R���n
��4�\D�(�zٻ�������9A����0[һL�4
_��S4���|H�GM_�V�?8q\�����_�<}'��f���-�USAx�n��)Z,��U���ćs{���{�u����(��StX	���9_	��E�wrzJa!fJ��Xu���;G�2|:�y}?R��oZ$Z��㣫���L~Ż�c�����HW*�W��Ed�M0��))��������[a��ԟD~;ZJ[�
�+�����2z!#>�࿲q[�1��5����gLyT\����P?g��מ���,`��4�_	�)������s������˭�,oQ�H�,h��0VRU<�tH4y^!�+5?�D��dY~�P�s��ԣ��z3�.߇� gZ}����OZ�UF�'?�#7�(%�!�򰨀D+�;`4C �v�� ���㸏��8��� `T�	�������ҧH?�t>���	?�~��������'2��[�h�[�՝���{����'DQ}�;j����<�����(&*��ߜ�ڑ]=��/,Y�6�١u�T4�(���Er%;����@1�P�sq4�d���#�x3��^���C@C��W���g��s���bG�7b2+�l ~��sU�țwJ=�(����i��2}��8>H�5�
��Im���e-���	�w1[U�
�A�� y��	]I @�v��eU@˙J�Ե��V����@ k>W���O�M�&2��L$!m��xj�yƗT&��T�}���W�a+��r�
b�@��a1����pβ��fO^�BN���d�*M��֩���',0~/Z��?�Vu�|�T��1綡`mȝ�-'����;�(�e��A2��ό�_��|w3U����Q��4���2��i�3�|���|!�(�b���!�Ѿ�T�ı��[��|%���Ni>�6���9�9�9�jg��`q��ǅA�_t�o�~���m�#f�T����Uȓ�d�2?���':o}P�6/~�� ��dfede$i ��Ct��^.���A�9���x��ύ��aܣ�
$�a���ț��r��"w�?/2�:��kadYΔM9Q����.UR)�\���g����;�&L�X��_w�����$�]��{�1�I���z���T3����#g3WMd�w�?;��D:�:pX̭t�8��v�L��<��� �4�%L;!��������,j��#1�EB1�Ox�h������J p?�e�]��(������fLl@�3���WQ���g�f�!c���d#-�x�>��G� UKEՓuץ8�_��;�2���L���om	�pQХ`yW$�?����0N�3*�B��'`�ѥ�,�<���N�W!�O�XT�s��iȹumf�49$�pb�#�������S�͇�D��Ԡ ���\Ww&�;��6�ƒ��e��z8���%�N^"���?̾���y;�Sz_Zߎ]�mJ-î�'����z��I�s���1(4|����#�6D�!l����=Q� qM��|�:0�K2����4��\�45g�s*^a=���.Xܪ��Y�^�^ne0sS���lbg�1f0�H��/��__�)U��4&��"�1M˟�.:G�����)p���Ⱡ!|���aP:d�z���cD-�wewK��Ѽ����������ۡ�=�6<��I������s���\g,�ZL���\ݫ��&��z�1l%�uMRu��M��: 0�@�Ӧ�M�W��D- 1/�<d{l��Ш�f��Y�Qu.�Y��V�2%#�OQ���O��D���|����� ������T�FNmM�_9cF��S�G����&T#�%cگ�J�\X.[N��}���,._������F)��_D0X�w������!�Κ�_E,o���\��y�<��q����d�iC";W�MhNvS��ч�r$?��:��?Ť��p�����Y�S�$�1+Q)�\�$��}7o����8�_������rO���˛u��]A�6Ϲ�I���N�h��xN��Րߏ�<����e�7$
��#��J�?�ʙ�O6Y�� CB��M��Q���r�_
SX+�CNl�%+$�W&��o🽗U��efO�&��0z"�GW�Ͼ�TX�P�,X�/��j��
q��5������/�U�Z���`�ݯ]��<��f��ƂT���˵$@�z`�N�����\^%�L���Ӗ���Pk�	_̙Bt �=~�}6�~�����+٤��Q��e���=��hj�.6�[���C����݆�^�8��C��k�M�=G�X�����߸�\�XN���#Q$Vm�
��Y��H�jl����P�����<*�k�sh��Dk��X�O�@�w_{}�U/)���".{��.�JW���E�chԅC����;��ۮ��Ԯ
�#L�I�-�P�XQ1��v��[�o�,e��(�Ni~��F�LYit�ѕ�߮���51�c/�M������'�V��[��N�s���걬~O��η��T���]q ��{�o��t�?��pLx7�n䐗N� �����:�_��j��T�|m�d'i�)�v�/�E��3��s�Jʫ�J
?���q����w�/93#λ/rɉ��D ���G��=Z��W�*�c)���Z�XHs�wwA��:��T���ް��6G�PzQG�q�C��������]wHk�L<ӄ7#F��a��#����0N1#��%�|��℠-	��LM��[�uq�g=���5�.���8���݉a��M��+C��,��j[�L���'�ĉ����
X��q�����oq%6BT�6�P�@�q���y��}���M���:S���R���`ij�в��&�|a� �����E�m��wJ��J8�n9[y��L����@ԡ�U
�5��)�[j;���>���V��4�1 	Xi�=�]��?��ܶY�a�9/;����,���lD�.�Dqa#63h�[�.��v��b�,�,�C�-
xF9�O�"v�A1<���_=*s� �B	�2��츂i�{§�D���՞�Y(f�h������R3j&�?Y�N���{�@�ܣ-Y��p1�)��w&�mfHcu��e:��T�����џ������|�������4}��)`7ϛ�$����:�}��~n.�Q��A�{r���/�5 ��>��{�I:��7%�C>�}7�2ɶ_劒�p�hu��A���M���<�zw�2�YM/ �<��;����7���8U$����?^m�x�:J�t���=H���\rZq7=�x�/K����!��V̓�k^���]+�2t��^�Xatx��Ja8��.9po�_��u_9v�h`c5��K�>r�eo:CN��H�5ݸ}�� �j�vq���qH4޻ֹD�b��|���S3��t�z%���0Q�~	=:�=����"��*��p���t���[�w�]�%����Z%N�#�f�~5e�@k����;&�"�l!���b�ƴ2Cd�s���u��^wr�r�rò�t�D:��6�eek7�]�;J�Y�ڷI �/Kf�^�����7�yr&�<I�{Ǐhv�JǗ�x��p��Đ��	{��֥ju�H=�.��杗�yD��N7X�a�E�a|��ԩD�c�k��VZ�K�;GK����e�8=$��M `2�'�4����`S�9�|Zy��E���W�Y��|Vg���_��2f���Z,�^��V���Jj������bc�')�`����X�J&��H��6�3r{a���'�/^�~�iq�ɀ=��j����F99G�P4U�?u�,��2F�ͪ�:uBt�	蚴G��:J�����^���ݟc�U��.S��#5���t��!ޯ�����n�~��[��B�\�P���$yS<R%��(j����|W�(�G��<v��X�F����t}�~�\ɚ�(����K��)�+�<��m��잝1(c�]<n��Fx��@�+��
�J^��=1��.���#��	��F�NA�(tg]�Dg�n~^���`f{K|�ZдdaBhC�d��`3U):�LS� �iԥׁ& !}���~�<��,��d PSL�p���]Yj��2�[�'
��.�-&����\̨��:�)�)C�{z��(�bF�~3�0��_?6!���7��$�GJa��D!�s���|j��='���#�����$���w#'�$Ph�:*]���ǀ�sǱ�3e~x��C%������C�xE�J:%�ɇ�N���O+#��v�"��H?n徝����W|���&`y6.Hh2�F��L:����1�3A��@H���-}�iv�@H��n���'Z�+�<�9	 p��b�6ݥ���F��)֧/ā�1X��g� � ���tl2y�{�i?{��ƍj����O�j��(��B�p��T,����΅WI�o�w��W�<�N5	y��5�#�3#�r!A�'ֶ���0��=d;����e͈���{u2���L�u%s)�(�{a�7,F�u7d��!6�~u䐴���0/��Ab���8P�%&I(gY&с_���bY�ድz
{L_G���L�b��{���b;�9�M��_I�^�?�h��,ץ\3F��m��l���Q��0�����V�~��[���aX����Qs!�k�Ng�͖�H�*:���V�7�+�1�Ӱo�9_�S��#j���v߽��ǭ�#�wdW� ޡ���TK���.o�^�X�ȼ(��V����3 ��~�8&�Է��q�}t�L����}�w &Ȁ�\���g�a����B~yO�jB�AU�08��N�/Ӷ���K{���c�"վ%�9���?��a��T�/������X������A��.x������Ɋ2�X�Q�+�fM%��^ ����EY�-��ln̻�ۓ�~���}���.�Zу|���'4T$w��aɈn���A<w5��"'�ٙd��h�B̻��5OJ�=� ���t���� 5�ﴩ���ʙ��A*I	���d��?H���(���G���າ��9V�������f��I�P�"�[v�|i��^nʂZb�5WG��m�S���x�]p5�M�[F ��w���՗Q=����+�H|q���[�!?�j�'�UF.ڔE�^�MynF�;�dE1��-��f`�}1�c�;�-^w"�����\��
���y��d[]����
�֡�^���������t�����g�v��q�"_-����9���ӯ�G�L���r+�_�;)l�5�a���c���π���$�z��݆iI��Zvɷ��@e���:�t��) Uz�2�� I�r
���z��$�L*�s��d7s8�6~�v�J�S�l�å��tzd3��wɖ�b	�v�%"�?n"����Kȏ,V����1��&�L{�m� g��x-A��	J�R�Ah�+�[K��Cak��.�Wg](���l=ΧiCs�8g��w�_�+�(Y����?��0:fܟ^O�nf�E��pB~�LYH�|5q��gJ��_�A��d�)a7�}Վ���z�xWͱ4U��2��?zը��\m���3�"�<�^A���/kU��������,���lJU� �Di��en[�`?��քv��#&�V��:�C���b��)=�z����`9|�q������Б�;
s���2YZ%|������m0���C�z��Za�����l/p �҇Y�'�\햒{)�8�jf�h�?g��_ٯ�B/�ϡg����󸃃*�y_�F�uR�IsL)~��6XZ������骪S��7����� ��T���r��^q5�ˏe�W�%+HmvJ���^�П�E���XO"���d���Qܐ�d�2�O����ɭC2�2j���9B� JX�n_W��Q��d'���5��ϰ�Ej����YH=%y�@
�0a��`�sG.��ҿ���Ĥ�k�w	�B7�R̛c���HƝ]� �`�k|�|)��͕A�)$�k �_��ޯD��wa�g��Rr)��q��K^}U��tp�����L���b�����]��Ì��S����K;
�]���U,�������|~���veX��#[��@&ol�1+��떚��'���52��@!�|���)]�(�95 ��U���#1urH��-��>\UxJ-�~�(�i���h���YE#w��{*�{�c�s�x��X6K�H�QS:�p��4��OT�m�TW�ɝ��Q��/���w~�(�����0�r�s� �|�τ�[P_/�D�,��;��3���b(�</�S�i�19�2��;��)��o%�&��-����t��s��6U����SJ6�F�J��o���\�#�B�z&�	��$AL �g�����<����[F�I�&��}�M�W��Q`�W�y[J�B]����c���OÅ�A���Q4�h�(��,�(�s��>�>!|YqM��9E����t��H��x}�)i��9?�9�����D�餃S$�R��tΙ�m�T	1�=�$p%�݌�TmC)l��8�v-Ù�v�.>�MeaD����,�*JDs�p��$[p�3�."�奔�:�$�2a��򲆋�{���6f�"��1���};�뤮w�&ܿj��`Zx�Yv�MC/=�C��u����L�R=_)&1�#�?���=#a/fj�~��&��[FrQ*2�����B�Y>n� è\�C��^�X$Sa���q��\�z.�U���(V��\�zDqt�IpY��2m�|�x��V���X2w��l�T��/�c���*��)�1���$ �{��Bg��.^8�Xz�@�Fw
Ǽ���`�	2$%J�®�2��q�s��D���6�7ɼ��<֞�"g��^�D��u�v ����8/Ñ�#A�w.�r���c�`/(��a�ɚ�ƭ&��� 4��������9���rp�0[�,)>�]H��s+�Ni�t�)'�蔅��j���|����*v*�#�5����;V򍄆���]~u:xy�{�s1�h���d`�-�a�Ok�~@�+[6^��|���(�����ok�^�6;t>Ȇ��phS�����%���%IEXEƷ�+|E+�[&��1�"��ֲ!à��P�=�[Tva-8����p��J���� )���|�kt��Q݋�Z
��x6�1C}f+E
	]�{r�c8ڼ���v��-�Wq�֛� �1ܱE�� �1���*h��^M�KAa���5=��][C;��v:;9%�SwY���:�x��a�0�ފ=L*g2�1��+�������]hW��PHYu����[�n�W�m
�T4&�	N|�/����j\�`��$�նT
��W�~��}԰�#4�4��b>g����~��}H���a��������Y�q{���au�B4B,�Cx���@ь�y,W5 N�w/}pX$���He���y���ƫ�"?�x��)���y�=q�����q|��^r����HXV�n%*�����;Y��P�ֲ��K�@:�J>�#��� �L�W��ԗ��h�S�|��S:�L����,�ζ�*��Oy)Q΢NŖQ.�*!�׊m?r1��]MP��)4[P���.Y%G�V����N�I��Y'U;Q����i��Ϛ9�;�ho�1�,f_�wP/��b�gI�Wj�4 �#�p;2�T2��<�AAW�h[r�O�������M0�`���9��R!�D�FÚ50�PNv��ȕor�d4J��Q+Ġ����|�)W�ds�/��VI쮭���$����x�?=S�M �w������U�ð2� K�ZA{o�j���K'L��&��9u�I���ӭ�����{�N
O�cD2G<��f�k<�w�1S�r�!�%KD�	络#� m�C��!��>���ܳ��Җ,�����V
�.JXk+;�vĀ��`F����)iA�w��ݩM~�A��K�'�X(�HUB��%�ݝ�(vV��It�GC�`��]����.�D�'�o�10�=���ң�FZ����l�G����w?��)���d�%�+��3g[�(�C Fp�=�d�O;U�w� v�3��jiۈ�B(.09���N�Ny��	�35�${%��8&�Gx�X_�S��+�y�#ZLj��N ��E�zj���bi��MW�}��xv�8���
�3}G]�(ڎ�¯���N��Bt����lw5��߉!�9<��W���x�@��?�l�ipU��[Sd��y��3�N�DM2���ݮ�/�c��2Y�)M�udl��l����VK����Pb��<͡~O?�X+fE�?�[h�bb�LX�j�ѲX�>)|w����a�u(�w�jXf�d%]�d_���tЦ{$��M�:�;z!KO�"�)Ǧ�Hmr�3��I���������Q1m?��9���� P��b>�:������u�@uUZ���h�L��*�)�h���E���������Ϙ�)M�GR��E� É5��C�����h�v�;CC���H�`ӿ��5�p4>�y�gER��"��܁��J\�uh��~�)D�Z"�E����[R\�D/����_&��H0�,��͊b����`�~��7t#V_f����ɜ���RՁ(�Ƨ`~��/F��uHж��_`�����Nq�o��ȯ¯v�!'�E$A��I*O�{TO=� X��Ʀn�!�AR`50�C $1��*�ɓ�O8��x��u�ϓ%n�j�(�,?�ƒ�V1|8�y/{���x��i���/���&N�Y�9h��#R�E���M�I�o�+<��'��n6"��E�WkDT�n�xo���@z�=�^�D�I]���&�Q�G\�����m�.b�p������3�fK
n���H��6F���.0����ӈ���~WQ#�{##n%���5-���9"�2VHV�ZxÀ3r�f#3��� ���i���K���d��Z7���n�Z��]��_���o����-[�[�N0;�}�[Y��"���N�m��t��d}5��p�6�t���Pzw�PMXz�fX%�+�T��d�f��͇H��F맔 #bD�(�!�@�ꝋ����s�KA:�˛���&�ҏNH����l����y8,�c~/�o����p���p�]�0F�5� ��$z�=��h�{��^"��^bD�6���^�ޑ�y��~�3��5k���\����}��=h[O5��!����)&L���F��ق(#�^�m�~;8��4fo�=�m
�����(g��9ē�{�q(uI)�pv2�H�喿QpO�{b7�6t���*�Q$�N�F�=������J��2&���s"�D�D-�ZO�w��Ivވ�4��?*��Ʌpb36��L���i��d9��_8��<�����1�>?��F2vy��$�EM����G�~n4
Y�G��ㄎgZ�26�B�sR~��v�����W+E1ubģ��Ru5LB%r��?�L��s�K��B���4�\	_*+MF1�+ik�ʍ�Ï��z=7����UIIoL:����h�m��'�����
�La]���9ON
l+ӓ1gE��z�-�O9ћ/^(i$��ώ1�v�ᶍ��g�W��w��q�L
����3��͝�M�lG�:o�{c��PP�u�F�2q#� 
��c+{s[����Jv=�(s��r�m�ZsSoF���C�d�f�g�a�SS#�+�Q2�^�x7D`�C�sѢp����|���n���̏���,ϡ�g}��O\�7��#�]`�ezl�*A���kGկ�G�UQ&���p��7P�y0N���un�8���$��+	���(��g��B�%��+�aͩ+(z���A�!b:���3�>�_Wj��9�a��ond��W�9G(	`G��N`���&]��]�<���K&ݘrq+t�ց�����t���}]��VU6ϻ����!ם������{��������\���W.d�������p@G�68�z�ԇ�.��ʀJ���pu��~����j x�Ѹi�m�"����JN�!;�����kX��uv^�}�eL�h��Y�����o���=���Yᪿ����g�\_�i����գ��R��4�LH����g�Z�S=ހ��_L<G^�;���Ŀ��M��A5��������k��H�	+t�1�xD��R�EhS�f0#�U
{�0�������	(��c=���ޟNW��k=nAG����>q�x�q��n>ZC-W��RqDvS��YC�-�	9(��+��S6�� '2P��s�q���6�����o�iY懟SGH�;R���V���S�Ad�O�" Z@(�І��'s#�	��0 �hR� �ˑJ ��;y�é�J�� ��r� _���;�gFF��2�����s��.[�,�8}J�8r�q`��X��/��y�
ϛ\�O_�|sk
2��sU���Ǔ��:7_�b����Z��QQJ��"���mb�|Ґ� og�����bq`��Oh��HGF����h/��q�2��/���z/\,Y������6 :$�� U���|`�Z7���g0��:�����)`A�"��u��Hq�x_��t1~�����9��?�8��.�E�����k�s�5�Oj���8|l���a���	�y�f��r�3����u�2]���L�r�1���T��i�,�a��aD
c��%��N-�.�\x�-�d���k��z�SX�m���w:QZ��L���>K}�{���ص:שRۏz�pՍ���(�����"��0&�0�@�!Dn�(�������ve��a*my����0H(a�#B�g��٘O��QF��O��㻼��a0����s�W~jf�T[���xɻ���w�o���|C������6���(A\3-��i�_
��5៉POs��%
���C�H�; h�����=�n3(��k�> ��b8z��F���P�����	͏�?��sMF����6�:Z�J�t���G1��e�*x$җ�-a�/~e�db����ڧ��g_|�m�o'����}�t8�?� W�$�Ec��i���*s�
��y��(`|��M�I��������#�n�M�j��u=o[�$���o�oJt�g����G��}6���7
�_�{%V�QY�2�̏�0�@:I	��Rg���i����0"�b�,�Q�L uz��jp�J"wy�R��#��r�E�`�:3N��f���V�3v��"��c	�S�z�J���=��@a�j�*��U2�������b�"����q��@��N|�@�4�Ժ`�n*^�.�sg�<�:�%7�Iҳ��]Ӝ" (��}ܻ�׆��a�}�T�1���v݁C,����{�����R�����qPt<��TB�t�B��޼���K���G���mV��*�ظց�'.�}b����"m���܋��⸤#�����wP��Տ�����x\y_;'='�b�M�9)�p=O��O��)�zg�1�]ߣ.���G�G�e��	6<f�$�\����V�5��;q`�����u�kOO�}���Y�Y���'Q��@y��D۴O%V)no�D]'t�
.!Z]�k*i^ҹ?H^E]�%��~i��R,D�/^��ʋsa������h�l�O�)���M  ��Q}�N3��)/���veJ6Dl:U���+����f�51��}P�"ق�>�)x?F#��ss�`k��W�+�|�'?ȑ���7�C�]�ZH�mP��ۺs7�E�#�f�<m�9#��ޖEZ'�ke�R�Ru��<],:���V� N<����>����x��MbK�Љ,�~��]�|b�fg2�LC.�]�O<bw�Ra���V�N������i��&���^����*U��p�:�Kz˝.���葥^k�4�={--�g���5��'yqq`�9�� ��_Gϑ���Gz�ء�c����V��0�����]���ݗ��W�sV�����&Qwt����v�9x+�+g6	L�>݈�v�ra��~�����a���l&���~�a�3�!��[ȯ���5���蚃��&�7�DPŒ��N>����3������a�.`�Ԗo��c�ZE�v���	�̧n�Nrzb0���z=��G����c���<��X`�q�$���|��^�7���Dw�D�!)!��RMeuV�?|Z��É��k�{z����y�V&���Zǔ�������!��Xo>��I��#��3e�?�*�yD\:J������w
w�L1mӑ*���`!��8nq]����W��b���3�AD���GNO���w�N�e�9~V|��(����i�$��]p3Zĵ��6�nJt^hg��_����}2��:�kax��]>o�A+���L�{ݐ؉ʭ�*��Q`��oU�5�h�3~M+ <���{Y��'���I�����`���
�	��/^���jb"[����}P�)vz
��ZxSo�j�`�y��+����8l��b��ow�Q'�Z�3�ʅ
�G�A�}���?pʪ����շk��"m�T�:X�ka�Jæ�K����'�36`��JZy��CL��=�	>j�*������4
m�6�W2�?���t)�0P�ᆳ0��6��O�	�>��o�Z�v�ޯ����W��~�8�|�������YL���Ť���^l�?`�`�g7���>�q�X�闡7�tS֙�`CD�߼�hUH�i]�J]�E��@�J�Y�ҩ���C];4�l�>��/y��=��խ���f����Ǟ�Ԇ�3;��a���E�k�5Y3�E��}\ŗ9t�b<�|l7��>|9�s����4T�_{K�6׍z<y��ȯn⹮�ds���jv璨J��by�<��j��}@ټ�N�������vaa\����:m�oH����Qx �i�p۷��.g**���S���U�A�382�&,��� N��l��L���[-�ƌ����)�A��7¾�EzE?�w�/Vw�E�(��TZ$�s^��C�Z'�@X����bK�1��r��8����������'Z�;�������.͈E׌bIA���RF��M#�d�D��M�*�$���x>��pP�G�`�
f͏��X��0�J8��<�ª-���:�s	/0?��%}��;����&��r��]U�.��Շ��&�Q%�Y1����u٩,���60E^�a���7a�\��|��lw]X��`�}��S]�c��Coȣ��j�z��8�a������������y^��(����6c�a�_��ӧ_��G�	�G�a�ja��X�҉z�ھ���yF$�fwl�+�?����۾����S����8��̑]��"-6	*P�Ԟ�}%�e���
km���Q�hW�L�=�+hY�#y�+�L��ꓛ��8C��O$OG�8 j�B��m����BZ]��1����:����*V�.�~�84��/j��>����7��?=4=\�P$��>#"��A-	$,Nnޟ3m�-_;�<Z�Z�z�p�F�t�K.�iM�:��-�ʽ:����RZo�loQ�Y�@>@t��h���%�w��w��j�|�\DX�Q%̮�Y�)C�ө�=�̪�aK�ʎ�N���7D־䨨0��z�	��M����o���\�z~�0����LGp
T�O{Ź�Et���92���Y���A�,s���R��4FK��������hk8�G}��n�T���(���4M&!_s�sɵ�8���h��U��;��{67��+|~����|�Ur͞`�d��[9h��_�˫
L����}�b�~Yf	LT��]e?T:������Z�]`Q���(��Y8��ݞ��G{N��@�� �5��O�>���[�����[T�{]���^&�r<�d"����z̼V�C�(�,�������8�k@��x�R߅�f=�8�r�b'���N�$��k��sH��;�ԞL�)2]|E�3��6�(aQ�c���OG 7��]h����B���{l�ׁ�j[�����|��[1�:�0�QlK^��us콼��4��K��,ţ1\tsvx��O�����:����%7�����
#&��j�E�dm6GW�4B���A�S�ϲO�yt�k幭Â�� A��aE��H�Bq!(�*1�V�o#�4&}q�b6ȔE �Lb�,�l����&���h5�_0�I�&�ソ
-o��n��L8�
�Է$v~^���ٯS�w�'�-�MyD4�:�b|
Ž���OƸ19t^{�ɸl����]t>�7�#v]-�?�N,Rp�Ƹp˴=�U���k��<D��͑Q����ĻG�	2f�F)`�)L�Su�og��2M\�=#�p��Z�\u�;�)����)�,�w���������Ny�	��~$G�o*s��%,����EU�qw��e�����Ҩ~v�އ��O�SM�Yq�Cǌ�*{�+�}��mB8��H��i�� �,��Ȳ��B��@�g6^��T1���Tϊщ#;�]I��66=�T�>=�o/ðxЙ�
W��\I�y|�aLr�4�1� �Bv1�g[蝹�Z�jm���V��[�C�I�ݱ�+�u��{a���-R���U%Ք���ub�<�'-M��xxʒ������ �}Y��n���y�W��	y�����@!w��o�୬��Ɵ��hR����]��B����.��
�pƅ.G���F�r��K}L«�z}�����Q�m F���FO���p���4���U���z洴Y_��.��'�(;����Ld�+n�I���>m�5�3U�����M�!D�g����MOo@k���|��0M�eZcq܎y����Rh�6tu���5^]��@g1�5~:����j���)4r�U���C��O2*���؞io4d���/�����;���C�\����f^�?�
��/�s���A���E��Y�%+Hd���g�\�Pvtj��b���_LM�?�u�Ӌ�;'��W���L݄���3��K@��A7\8�ߨ.MBM��oV��n%��*ͺ.5��CKL\kLk�Vq��x��=V�T��s�E�b�qڶ�2YxzU�Dp+Ir�K�p۶7Hʭ��F̘�i���r�E��z��N�XxO�����ໞxA�l�/
Lܣޕ��"��Li�=�*��ܯ_�j�vK��Vԝ�Ye��f���<�'{^�.nܐ��xK۸�����a�N��lb/������ªWc���:��P��y�ΓXM�*Ƭ@��fX-�Ա��#�������-�
J�9�)╋e��ZA�Oc�{�､L�Y�۹�b��Yw�x_O���hv��QE��"tN��\��{�S�Q��E!hj�g\_r���cE���|�v*�f��"V;��+����&#-q�}��p��%����6�#d��GU4LJqT���#�뛗 ���oۑa�A��ٮ��!�.��2�w��m�2�I7��;��s~�2�^�?  ;�5�E|���˟ܰ:�V;�$˴ly�|�͏�or͇0lo�*	��bRD��NP��+�����*jE7`Z�.R5�&�.�N[F,���)OX]�D�O��e�E��D�=�Ǝk����#���:xl�9�D}�)x4����$��������b ݖ����]���f��bx�VB�5I�pV3�7�r�I�؝���O�6iY�֥�R]�y����S0K��?4!N����l�Qw�=8i`(��{�(�~w{�]�zt�[ A�����g���MX�|���Iviw�=���hG��J�'���c^��~j}���Jr�h��I8�g�2m�{���J�I��b'�˯�C�_���*��1js�zCS��Yv8[�		viKL
��~�!�h_�Қ��0_�Dxw�\%��
�T~*ڎ�u=��MB�czC͟�٣��5m��8�y�5�苛��n�en6�Q��FG	��;��"����k�	�)��(w,�%�F�Io�k8��Q�jr��ar����;~��!�##>*�.���0�{�<zuKf�ˤ�B��q��	�x#�,��'L�m	�����ti�Y�~�B�:�7y���ǸY7N/^�=r>ZC3_�K�o���H�!>l!��,�^�ȍ�-Wi��;�Sm�mچ)ԧ��3
>��i⧧��d=�#�wΣ��KB^�R7�f�ti[.s�Jv���Zd�p���m+is�9Z`��%A{b��S�k��v_��<-�I/q����E�H�Pȥ8���y��#V�܄.�U�v���P=�\Z�O20|�m�^|��QR� �qع�mh[���i���;r��oׇ�dfGr�t�����z�3���:t�;�FZ�&��6�:^G��X�"�����M��3���r�[�����덫��ʏ�2�c�Q!.��Ac�����o���Ez��}j�w]ƚ W���Y�SZ(����\R�:��b��vymÊ@����tfr���$_;>���۱E8�nbrxZ�G;�xZc!�����t#����ƖT%�M!����h�.9�u�{~��z"֫���j��%\�;.�F��ZE�~��V��8��s�C� pDk�2��\���@6��豱����Nr1᧗}�@�qQ��~�|uay6�(�_���K���*��~��{;�S�Է �z�y��"��l�9+>�X�JW��'�dh�⑈���O	��ܯ�i+��T�E�Q��gex;X�Q��G��_I�ӧ�T��w��EmZ+�{�^�5֐D��g���1�1vg/iv��PiH#?L�ܟ�N�W�7�Ė7�Md1j��rU�������a.�~���dfn�U�d>����\�.u�^�N��QW��u�-,��dɿ���
%��?�_}�?^�qոsQ٠�l#�q@8x>Ї�]
�uJ�O{7���g�n�P�|�h�z���#��-��U��t�3sw�����g_��6�5�`|Kib�i��������L�F,�b-��6��}'�����8:$m�X��_�eɘ �B���R.�
�&���w��;�3�I���z9#�8U�DƟ�Ѥ<�.T�0���M�o{��I������L0M8 ���ɷ?���\@���ig�5��c�hq���o��}�$g/T�Fĳ|�p�<��pu���Sn�Օ
�jA�V��&Y�]U�J1�Q.��nD�d&�f���H�l���A/����.Y~�6�u�^9��F':�=1ɖ�)�}ˊ�����C�\:�o+`Aly�L%��%*���t1�i4���5X}�T�S�e@�I�O�u��R��֙s����p�` WW�]M�#|@M�������Mv@�HxO�S+����*Ł�֢�w�G�Ɖ��<��p쑼�%�t�޿9)�o�c���Z��K%Ya]�בp��������K�6%r��~�� �}	���G|�C=��3�>_��ßcQ	��ׄl��J~��h�V ��h3J���k%�لuTxqv���Bʁ9��w0�t�h�A��1�~Q1��'��L�[˘z���="�.�$�nd�`D��E�o��gF���4�?dXߵ�KR�B�\E�g��7LU�_��ƅ��n�"�N��Z�$-��6�؇��D�(�|�Xn��03���fX��nc�|�'3�5���e�f��F��9��:��]�Vd�F;�KI���v���#�,W�D�?��{d��$�
�Ѻ���S�Y��E��.���՛�a���h�Yy` �uE17rHxf�9���v´�͌��~�&��6K���r����g|����3wZ��М��q^%�%gS�먀2DAH4����V*W�n����$�$������(��j�y"�F�;�h�\�@_�G$�^����Cn�gm��mؼy��1Fjצ�z�i�G<���(���ށJ+�D��L5��1��h	Ǭ0ͮ3����74��Г~]f��Z�^����-z��:��ρuY{e��׊�#u�W6.��	<Ru��rv�E��^�u�ԅ�t��K�fT"�=D�|�|(66�]=d��[3T�еoĺ��o@�kKu`�]�X�uJ-�H�~���=?��X�K�z�E���A�,��/��*r��Ն��2{p��XzB��g;W�F�^��(��FU�e������[�QƭQh.im8E���"����s��jGA>�RxND�P��vO�>���
1��W��~3e����U��.T}l�PW+��vT6\v�$5�`�0���Ɉx�t�4ʈ��9���}靊::�D!��C�������Y�:U�XI�ϊ�J0��D[�!�	��𪾉D���M��J��F����m��d�k"��:.'3k��Ñ���]��xb�>����/GM��ӿ�@����L
�ߤ�VA�ɡ[�;��A!Z�&�#k�u �)�b��z�6�X0{�Z���:ꠙGFK�q9F��Nڭr�9=yD"�!���C���/~���S�=J�\aJ|+A�T[3m��2\/Ǣ�S:;���-��Gǋ�.�߹�$b��۵��h ���=�}�'�_��(�U]WwO��7B�_�^2ʋ:�m��uB�Ǐ�R�8�Di@.����۶X}=��q}���ø�ϨGP7���|f�^��?{�q8���WX��{3�Ʋ�d������B�E h�#�>�xKQn��rJ�J�6`w�.
�Z�V�q>��0����Beru�K���Q�o�.>�z�AH�p����C���/*ÇOָ?��罗.����ov�������˰��ܽ� �����*����IF[�Q��˥�B�/8)~���.[� ���
fBTn�W�`����Z����l9T��hN��	̃5uwh�()�[sꊢ�I(Z�b�wi������?i]�߬�����c$UO~U�	2lEadr���h%��pv�㱕�|��������S|Ҹñ@�-d]��Ux�M��3��'�:etp��\|�+�~+�![����	�<r�h��Tf1�WS�n�<���
e�d���vE�m�G�T}�U�ox�9�C2�;�%������g�Q2����A�!{�o2���P<����^�pW9cr�$˄ %�nډx9���U��P�L5��W(��k�C�2'�1�4^��r�hJ�a�k7�

��~�S7J���)��F9��B�l��ʉr�^��ֻ�hj0��M���s�)��5��cM'6�"� l�c��c��tͷCM�$d}��� ]$������~�_�z�]AzW�@P�J2C!w���^�m
i`�"��?�� }� �=;���t]s`����;����1��-+�����12�Q[����H����uzX��_�~�_��!��h� ��LUw�5�)����C�,s:���֫N,L{��@!�f!v}F$0���[C�����F�r���Ͻ�a�|7������;u^��A}VY��Rï����Ff�u�sirj�s����Gn�O,9��r&�Q0��(>�<�ną~j�uO�q괘�'i6u2�-ߖ�w�")�h�׹i����d}�:�߲,󓇤�gh����� ;�'�h��ium�R� *�9���ۤ��d �U��4�����Ǩ��/Ds9����jN�I �>UGG3U��X��'b2m�eܝ���:$�R��V��0� ��ܒ�&�,y0����g�Pת�@)����!r����_�7��:wr��L��pa�����2��׊}�C����P8��ŤQƩ7˘:wF�=� F��i�����Gݹu5��ӫ�2Q<w�U����1���k��J�4?�'@P�Љ�o��	J���[�����E*�
��%�<1����}�Ł�x���?��~]� u�����@ܧ��{/�^3qǱ�e�Hr�\9n��d��
��E�}<\��`*�vAx������q]��,�%`A�,�2f���(��8�Ϸ�D����ı�ȫ~~�!B���<�4O��N����,�=�q�A� z_��]������*�$��P�*��?L��\K)������:6����/��: �A���[$����I
6p��ڏ_�W^����c3���{��r�ev���#�	x�F�SQ�)O!�/;|�s�OQ�_��<h�$�Kk #: wc��2������ϕ\	��F>X��ש��� j�HN���.��8�-x���0������
�`�߮�������wYڄ�3 OlZ�h�� 4Y��$<�")��74��'�ٳ��>�Gh��7|���S�<[u���Ϲ�a�塇��{\-ӵ)���t��w�oZ�{��Hʉ�����x�����#�]Ʌ��*X�CeL���_��f�c}";�ȧXb���R1��xF=�Sr�5�)0!WH�r� =�������.���t��������3Du�����v��d��È^Bx�Z^�P/nj*c��ݗ(it�NxQ���5g&��3�m�K)�T�ǉ�"��AZ�"�؁��;�t��A^�~�r���Kba�%�� �d�~y�㹊	��Z�qOSlYfz6�BwSQ�����<��͏�AjqQ�B�4'i��6��\��K3�������pzT�lI����A�L���Ր��-��\�Փ5%�Z�HHXb�J�������##Ξ���{;>�<�}9�0 �s�����<pý���ǹ%5� �ђ�օ��~dn�s�E� �,b��vt5�i ���^xf�S���N��Tn�[r�e�	�9<� ���%��|F�gH�6{��IM��7/VY�&�+��C?��d��e�8R�o��=�$�l�4b03���R��fB���0�H0 j=�;��4��s�ʞ�71X(>#rː�����-�ԧo�ר�%^D<E�x��"H�GL]Zp@	1�T(ВN��7��*��o|��@����l��{E��S�T�<(-bC`E�g��W�߇�9~�ߊȱ�.�^�9�|��Ɲ~w�"ȆL���ׄ�r!G�5��>��%�+�vcʹ�Gc�W�6(E3|�up������Nէ3�3G2��ϼ�%��3���r2�������؊C<J�1�$-����D�ݭW9�ƟH�v���Om�
���E0?-%ӾPc�*�;��+*A�'��R���z��܉WSAT?S02����0��%b����ޛj�5�48}�^�}y0��B*�P�k"8�*�^���ԥ��q�î�e�´������ԝ��џ�Xik�5M�G-��^��=Q�WWta��*�ކml�/e۽Y�vtz����=�Q�_I︵|���q=r�'Wy5ɬ`F�C���O@�p���A���|�.!��<f��8�-A�����X)�8D(���}|�}������vVt� }��4��	Em6,�Q�KJT���(�y��]]�-�#L���r�ź�Q��T�L��A�0���X�k���p
ק��o|���ˢTg��1�Q鋏b�Đ��Gw�����F�^��$�M�1M<�ys��"(A8΃��U��>����k���ڡ74f���xٸ�w)P���=��˙�S�'��gt-PO��"�ȉ_�*b����^�������zL� z�Y�M]�3�&u�w��Y��eSL#��]�����,&���3���oZ���+\����_�~��J�2�:��~P7p�S7�	�֤:$b��Um�P�Fg#W�/2�FD�蕷��e�����4f��=�f��qZ�]����'���۲LvQ}JH���[BR;�ņ���[@о����xHǒ[�������(7ޣi��\E��{�TU�^^H ﮐ�=L�wL�|%���7�|�h��<Ba��<sx�OK$0T�:��co��]ޗ�|�U�l�����ͱ������G��ը�~rF3��y�M1߰�lƐ ���7n����T�+���u�h2�~;�R��2�����^��d6��݋N|��#�snJ���kE��tk�-�e�C�9C�J5�]W�(�oT�S�'�����zN��%�GAtl-�4��P�:aNp�ܾ��� [=�y0=������qR1D}m���iY�0�Úb�Et�$��K�`K�uB�hm��B���0*��2�=Oɗ��ƨX�B�-h	=�K�~t��\�^�S�<B����mW���Q�(�m6[!kk����GF	��=Xq�L�#���;�D�mS���f��M�z0(am�xY�}��~�bQ���M�ݒ2�ÿ������ή�ݥOR5KQ��^��������@����i(�=��������m�C'*��ؤt��?ḧ́nMI^HK�@�U)�r0�Y�� ��Ɛ�k4.����O���U��4*�{�7j �����9��O/EP,�ΥW���ϣ�]:H�+��Z�m�Lo�Igd�r�K>�r�jUW4_,(�}��4u~J��xuo��l�#PP�L�J��k�@U@����X>�:����3O�[�a樼a�e���'@1:���*U�U��hrVvF��9_���S2�N�`�/�\�%�[�7�Zg�P9��vd��.zm�dՓ�ND��,�|;�����%z���8�p.~���ܟ>��U�u{~���Uw�@xG���ֳ6ɒ	q�pWn�U��<�^���n9[%���rtS��	�����Nt'=�4_�H ��D����D�F���U޿oZ�K��<�gY�A 9n'~B]|�@<�?�>�{�ي�Ty`<8��-�bus��K�uԫ�m�C<�eD96?١^��y瓹x��ɥ\��{��נz��,�vL.>c��?��-t��4�%V;|�~�����6]�z!�Ϡ*D+:q�/`�1�M��Ğ�Ѵ^hJ&�߆���)}�:�>�������R�?o<Q�̏>x�n�>D�Ln�����ߑ�MW�i��N.r�D��<9�+�B{��Q|yЧ����c�����@RV���hZ{F|e��꼗�F�a����ծ���䃐�L2FF츑�o��)����m/>�+U�C¶�nW��,-�S�M�Mpў���@=��X��<Z�����4ݎ;��}���f[��ʗ���C���J�R��v>�1�	|"�j����d�����d�N��̕.����W����^�E72H8>ɪ�doT�������aj�F��*B�F���)��n���O�+�x���������d��Ղ�q���EA����9۽B2���B+|E�)�c
"0��8y���|��<�>o�� 蘚{�h�>� ���tS�fU汙�\�7{�_;�R�\]d@q�Et�����N�K�� �(y�#� ���+9��z��/�4�:��ڪ-k�u]�9yxC]N���"���kh��F^my�L(i�UN�W��j�����/HD�/W��7�4�%
�_����;����gz徐-��\qA|	2sV~�rdώ���^Uw��Z�K䢶�4�s��+��	��%�
�PϚ�%�r�F>��E�e �s���#����u�_e@s�D�?��{_��Z$z���ֿP?UV��Iu��Z��S�sY!�YZ+WNM-2��k*�vV%�I�o�-'0�Yw{s��E�oak%�O�Mw���P�W��Mf�����A�t��Z~�o����6=`��*`��"���v��'���L�G���Ѝ޹tҬ�@쿑�)�m?���m�uC�J�֟>�N�ѫ�����%^ۑAXA��'���3�����U`��"r�j)�)���`�8�G�r��=#ºa�R��������`-��A�;����݃k�����T@xc�S}��C�� �oQ:�~OW�<��� p��r�h#��=�<8��6��n��5W��&=�/>0�����2U�@!�r�I�ڟ?�LF�P�U��YUFg+�`��s�%C��<������O�y�Ӑ���sn�Li�����lTg�G� �fH���\E{d���=@�w�4~@�g+n�<���� �`�,����f��ߜ�h�*��aB�-�)��{L8L��h��x��tk� ��D����Nxl[�P������+�*���pr��d<���)�V\~�A�*+U�=趴���M�~͈�5��x8_�ڋ��e-�]��܌C/�f�Ws(��q�|h�������iaP��I--֮��/����Ga��q��!9�Y,�UR�d쑵�{e�܄x�������M狣��'CҼ������uH�j����kz����h�]��B�������m�7G������"� 7��kOjAWQj��&�[�S��&�i�!��4oE����m�M�)���B�0���L�ج�L����r���zno����y_;jKŐ���=�$��Za~p�s����ϗ�o�� m��}b���$��l]�}�N_�����=��B�<���0�>�f��m�=�.O����������	����u��?'՝��=8@$�����_E-ҩ?����7���� Ax���;�ې�N����AM̧laѵ�4����?�>q����޻���	�Xx�b~ǆ�;:�{��r!�>&9�����m�(#N�^Q���~��%D�tf�����zc]_�]u�MB��ٙ0�N*�*՞���Il7�����*c���ZA#��}^�GE%b�k��s��[�IWg��սI_��S*�e���Ќ�;��`U�qH�n�SCf:�{���u��0��	��D��%i�'���@�T�!܎��P�.�X���)�a�t���2ZP-!��{�)�`i��1�5�Nu�G��2Y�����lZ�jrGS� ���S��sNN��ߞ�10�mڳπ�	�����Q8���]���o�2i7�4R�G�썧IoSXChz`��3E�x�K'��b>㨯��S�@-w��G����$g���|"����~�U�?ן� OI��?ݝ�)�p'��bز�H��혦�<>�xm�� �pv�3raw�1rg}3��\��: U����{&����fY?3C|�������7I̞V�(�S�l��4e����x��ܟb��^��^��F�C�0s�%�$A�=�f�Uo@���ކDᝠ"���M�D^M�:�����U ȢC���띷�4�{�p�1tKk�!�Ϯ�����CGW�}R�ߝ�n�g#H��<K��9�$����ˌݖ�T�1�;�tM�k6��%�����5�"�5�k�MδZ��Z�ȏ�YO�r��>!��x��@M�L�Ʊ��»�"w*͹��n���ƈ��0z��W2��U�M�j����� J������\'ܭ���.��'"殯�s��;�G=}�4�w��{0�Z�;X�E�<�Tz\t��B'���<�����1�~m���F~t��Y2���_��TF{wb{*ж��Psh��;�q�:wm�];>p���U�B/�4�u���m˘U���*���%�k$v����h�-f�򭙲�������� �7ڨ��y����9�wZ`�Վ �>����6dt-#�*ɒꙨ�mr���lDhC�u=��뷨�&w���-�D���oa��>I>�Y�s��T��ʊ��p�cE�7"�l.��kh���S&-2*d�=O;���o�%���O㭲�	�Y{s;jίh�w%���w.���������Ϭ.?ai�� �3�d����,)@��d�5M@G$U��')5�'36��E�/c�*l��م�����tq��v>5C�iYr��4s># ���%�2%�>�� "oI�s������N�.{��T ���L�YNPb�Wi7Υ�	/r�/Vg��T��u}p�6�¯�P;�%����ϫ���c<�]�.ke\��0*�V��߿�W9�dL����g2�bW���ne��a���'�#&�}�(��	��yW�xy˰(�.lX@�F�������P�������CE��n�.���{?��=�������a�}ź�:�y��`t/^q�u7o6�R ��[�5G�����T}��}) ��>��F�/ܹ��;�p[��Q��\njL����攮����DX)Z*���栘}��,�ӊ�w�`����c`�����W�I-1N~W���;.K�^���׫Ɖ����o��,���K�bת>�,�!��1�I���ʍ1X�=����K�ꊃ�ŊE�����=��f6��r[_*�1�{�⃁������X:X��������Ƹ���D��1
���(u��*�vk~ݽ7����l��WhnV�1���t�mr˘eϢ<�J���lK�7����s�	j�K(z�W���ME^�@�l3���D�&wʛ�ʟ5��G#~���o2*-�tFվw��C5�N��H ���q��P���?�`,fd���0V�P�X�8�ۮ�,���Ms,��>T��V�����Zo�,<�R����c6/�hj�4�?�ۮ�am������v<�9���f�������{4�z�Y�7�O�S�mZ�LYUs���t�u?,�_��fU��ҟ��+��<��^_Ζ�&�>U���z2&x�V�#]��őAn9�k��l�Q��ID���O�@u�u&��r��(BK���q�E#�D~�#_�5�e+��G�i�5�1-}���e���V �6�0)Ilc!�g,�r����Шu����*�|A��+��b��:��z=� M	8�'-D~�w�ou�|Eԕ�F�w���vXj�����@2��F�(L_`K�y�/.g����8-�_�����j1��ZV��o1{�E�Պ|clɶh��������ymQ�#�@�����aq�[$�&p[�ڮ�?��"�L#�n�C~݋�#-�ŉ�ؚW���҃k�3ځ�`5��6(�,�b;�4t��u��q�����@,.���A�B.�d�V���%qΐ�W�y���ʆK�W�z8~�n����rFi˨n||����K^�+��@�����m��T�04�wab*�\u��DB�5�����*�x:��������"U��S�q,?�u~m!Z�5]T1ZO]l��C�ǻN�-6q���~6�+BP�b6v��d������ ġ�2Nĭ����r�6���~�d	0MQ����M3����d�
ͷ?��?_>|1)g�����G(�����[��T��T�[�Z���<�C�a�;�E_=�B��d�8�LaȁiY��f����;��"��pb�]�uF�����|g C���M�7N�ETb*mHnoJw�@�¥,"fH��_�`���?��nӂX�7��D��0��Tg����{���Z�i����W�/jRx��FttFIz�Y�1i���2��_�g�����P,SЁg�ZK�j�eH,B  �RES�F�ָ���ęu�V3��&���5�/�"d>InC��Ia��]M�q�M����YV�!q�o�O|*X�O�R��)Vr���Ԣ��gp�X9�u�g�����T��ls��T]�l�v�rv�])�FP������H)DmnN�]�o��=���&��U8�����M]}_���ꬱG>z
�>��a�J����Ջ��gާ�E���]����[lHFwލ ��\��ȇ�Vd�璧HY���T�=�FӪ�d�&�pӷ��]���^��ţ�W�_i�xJ�ST@�Z.w`���m�nQ{����=�&�@S�;�v�흯����;?V�c�&f�$U�:}�r��������ܝ1�ޮ��7G69�Aw�ޯ�G�g��1}���Ӷ�%�g����-��_S�����:j9�i	�P]�(��6�������~$�[ʆ��m)�	�����.�]���Ck�a?��22>�駅��jUi)Oq#� �4't�]�eú�a�Q�_��_��R�n���^�*!8N�H���ݒ�N*\t��x/�k|��/����?.8D��I������O�s�T���Qu����0�S��������h�~���q9
.9�
x�$�ΏGtzLؿN�a�J,N8�cZ���Q�ù^�Ǎ�A�Am�����Ms��t��Ĳ7X��>��Ȥ�;q�h֔���U�/J��N-j�W��v.`Ž�z�.�[y�q�E� !^���9*[���E�ڥ��A��ږ��`v��l�	�Ū�O���td�VH.���K���W�Zh��ӎMB�>sE%_��k|k�Ζ��N|#q�T��5����C�#͞���w���z�[�_%����/xG���_wZ�-&��k�G�_��3r!��~tKd���\<DC,6���jZ�I�)��*�\��[:�r���.M��_{<%��p4 �l݋����ʦ�5ހ���*�;|X��I�^�@/�|UZ�X�e��:X����1���Cx<^�T{�8��b��E�h<��ߜB�ie5����Ś4��W�~ "x�&��VZ�
�Ub�Ľ���k�Z���N�&_$�!g߇z� 4Z�}s�b6r�2�����u6w%�� ��r����P	Ss�L^�	1�K�B����i���-����?�%�FK�!���
Zk�7�DB��ڸؿm�6T�|v��*s������J�~�� }r�D�[���0��Q�?�g��R�F�t�#�9�#��b�r����zW���mD����q��N�.�M=�̪2i�˞��l9�ԯ���K�6�e!˒0��3��7�'���Ytw��;q�Hb���J	I(^~�Yr�3n $�R<n��؄9N׮�X�#��������X́a 4�;	rKk/E+`8��*�.y�+�n�Ǵ��� �/ge���������NhDUa7�S�zu�~i7K���#��6�5��\=� �i�jko��V����Q�s����
@�\WË�:��ώ�ޓ�.�-Xc1#�M��N|�z=Ū�Q�Eʎ_AW�0���^�S��ַ����5i�̣�Rě�e�%�����Hbn��5T�?G����j����ž\�n�����M|}��Tk���cN��Ye`�a⽗2��8	m��[=8�+��ީ��K���}�͖�Ic��;�0����pk3��y.L\/a�i-a���1u�e"�x�0�f�?���Tג�3a��a;���N�o�t���L�� # ����C=g����^����,MCs�V�j���/h��A�5��pQ����t��sg��D����Q���%-�l�pcT}w��%[[��ɓ��!Vul�	ժ���k�;~H�Γ�����VӚ�v�/1�~1��ū"б�Y�lV#�w�.D�p�N���l�կ29 R�z��,���K��͛��]�,V��RX-�/B�zLf���A5D���
�?qg����s���v�����_@Α�5��<�5+_�R�b�ؼ��='<.�_�5����ӃYG+=fK��!�a��"�.K� ��=�%�~ 꺦5І8�y(5�l�NTe`�m�LO[�����X�~6or�&=A�E�����J��b�[]�5l!��w�ַ�d߫����~o�i����F#>��\M�������{�����3�Ұ��^82���Jo���>]!M6��O�0�F����R+�������ycU�2�<�yb%�tQ)-I�
	�]���/���/S�E:��)�P�Nu�?��w�ü�]B�D�V:������i�7�ܓ���
���7@T>��7Ջ�J��N�od2I�d3=W��������=�5����qiw�\��)�6�Ի	( �oB��7s_e�Ǫ_��k�=Z�����+���q����<�1�k�Ԗ�P鶑=�(E�KW���*�_�#I'���s��<�eد[0��L�9�v�Ν����D�C�����D|��a�;w�%�~5��R�i",�/���~r���' g7�R�6�O�]�T���J��Y�v���b8W��f�FV��� �F��9�XTV��`�]�դE�r�SA�#��x�����|�k��'�_��3SL���A�߲��+���G��3՝.��_��d-�@C�K��AΗ�ǒ�%h��1w���{L�����7}�!GpƲ��K_��n�Ra��$����}G�Zj<��M��ʆ�{���-]+X��A���z��E&��2��9*ߺ�=���+s-<���e/�����[�[�١zWg�_T��%�%~�ó������ը��U3���J��ͅ�`�P]�K�s�/���W1ʜ�&�ͱ��Â�V\)�2�ە(N��>��^s.Z�"#����>�A�~׏�uy�ð��ǺK�izp�C���g��H�S�-q�B���>}�����%��;��&\�ѹ��������s�5F{}m��a��9�=O�eB/��:hX����h��2����ͼ�@���{��JCΜ}�ɮU`<�l�is�(7jB��0��>쯴�ף.b��G��hx�iSQ�y�2��]Hc(�����<��}�W{�׏�X�V����Q�# Q�K��+���$R\�
>�����~�H8<���z����mFe��p�[PK6���ܮ��u��T�����Z��y�Ocu�[S��/?�Mx�|�"u�iլR���="]�j�o��}�LgY%."�X�x���?զ@B�6��7�L�j~ĉ:�[l�`L	 J�ECK�5k�r��:�� ��b��p��2�|���i�/qǅ�Nb�	u&":��U?�3G?�Xϖ:��\���?`�/��Ns��1߳L��d�����\!�{���~�em3��1�*D��K簇��G�;���� ?0f=�Zڪ��W���o)K��������I�y1�_�>�^��0���M��f +Ծ��d�춣|��G�n�4#�|��ё���$]�:,��.��i��p3*5wu����%������j��g��p���'���/�%'l�����4���/-��Ѥ"��4{�g����?���=#M�3
���T���c��dw>��l]�m%Ud�����"��$_� ��`@�?�w��ȔM�23�4�H?/4�Q[l�<5ͥ�Z�T{�\n/��N�Y����\#�o�x�/�c8aL�D�&-�<MY}
$��n�*� �vG#�ߘ��OHvK�J�K�|���  s����Z�%@��+�+K�I�Y���O��v@�T<�O�]Ň~\��u3�'�Ȍ�@���
����4+/�@6(��J<m�����1�����L���v{������2sVY�1 ;�r���/�I������PecBAE��?y&�9�l&פ�$��}�A�v�[��ez<:����g~�Pǳ��`$}��h��Z�!U�C�1��<p�LBg%,xK�Ja����.��L�7���oG��-�bV��rR������`+]�94�l7��r B?'{�]Ws�Nt�ZiXҨ� 8���(@�d ��@����9z����Lm��<І�`�̓���a�H��]"X��E �EMo��s[#�:�Ў���P,t�'_��uؘ��9Y�p8�L9\��K}甫���8�����jn��t/�B����֖@��������m��r���d[�ds�pz������߭�JV��P'KVڍ+s�6J�cC���h'B,PI��~���J0t�T�c�8 �mɱ%fٍ&�I�r[&��m��A�rj5�9��k�<�*��i��L�ƅ�ym�X%���?����x���<�	ZD�_����z	�������Ȧ(m�g/u�{WBx�2K[�,��r��+Z�k���:]�|"b��{�"Ãц�an-�@e4fe
/�>H�=�B�[��=�pM��5G���d�#�ޗ�la�'[����O�9NqV?y~�uLm���hם����b�_�@�|43iY]]ny�P�4778��Q��ʼ�F�L$��aya�F��t�J[��y��S�*��XSM�9w���8q�zC�p�u����cTX���:kd���G��;�ڧ�����L�t��Ͽ2��M
HV�&�����Y3��*-���>\�i}�YW9]i����}��������y��b�Vz���NN��I��Q�u���������A��,�-���gīO�Y��>�y-q��m��d����9+�F��3�ϣ��'3�؆>aU����5�������`������
pKg�.\�[���	�d��x%�#P�Dd�.��������~��4��`����2iM�Ͳ��͐����/Lg����Eew��������ؚ�ݯ����l#XQ'�ϱ�<1� 	��FQB��V��ڏkϿ|�c�,�3^315���ѳȨ���
��: ��F]ju�.���_������p6r�FW�i�˼�1�Le�����~�l�b����C-�"߮��a$b�����g&��X9�<rϣ��̇�)ؑ�qj T��]`n�;=��~to���g��r;7�\�ꪰqve�Vb��5�������G������ll1ܚ�|���N�U������_ӥ���c+�FϫՎ�����c;�qc*Zje�h���eGQ�a��A뗢�}!��-�iB%W��]P��ņ`��,=��/�d�G��v/.3�ı�ݡ�\��fI���|�"rg,����[�C��\�q�p8l�S�M?'N�*���=�M`~�����u1 ��6>YY��]�=c��e������.W������9��o���0�S���Y��d�u�'&��~ݍѭńd�Gt,���{����]�8��Ǣ�ѓEүT�/�����~
'�y��Un\���45f�ɈC�56dKM��ؼޫ��U���2b�"�Sܭ.4�Ams츋Һ��9Pj������~��̊������<�����V�G���L[���%�=�95pD���㏼x|�A̩��<4��~��mQ�t z��S ����1�Q��~�|��y$�w�Oz��BQ���ǘ���`|0�$��R,��1�D"�W�	��欏0�*�ӨH����c���s��~�7zg���S8�6��U���҃!{���4r��mq����M��ݢ�-ڌ�I�?�f��w�G����$���������cY���
���J������?���q����S����`[!$�fO�� �� H=߽	橈~L�����?S�_�xe=�����p����!��c�No:�Kp�����Ά�n�m҃���N2���G`׫��`���m�a�_P�m�ϑ%���/�*�Ȇ/����@Dw_g��e�\d!�������z�s����?�B���x����S�Dt�~��v��i@��_YQ����	�U�VM����Ȯ�F��iW��f +\Gk]ᅋ��� :y\޴<�H����퐍7�a��l�����<Q&��{�� ��Y\gE� `���i}����t��W�����v��z��c���_UC�a�vu4k�I���P�o�"����!o��-R���z�W�?33O��>���q	/��lȚ��t�3�9::%|��:)�V;����<���ج�nc�!KX;M��<�j�&lr�����Ѣ˲���zT��>�L$�Na�U�pK��=|���8m�N��{��o�t��;k؋(�~�*����������"ecП�y�I�����r��Y���v�����ï��i��oM����ځ�S�ݓ�-WM�rc=�6�*	F�N�N�vQ#�=чs9E����=X|iʝ����x�-(�����}GG�ûo<�1����o~W�Fq�S�S,��ſ�@u$S<����-o�S��Ӎ�e]�,��,���Ag�aw�����'������|�[H��pIkjWc�5��ge����	���@��D���2�����p62��L﫣>����Qz�!Y��:����fk�����M�4�����,�Wi�͔�\��6	��x�c0�-Z�@��!0�@�cT��Lb�ٽ����^���"}���RvA0�g�t(I�z=�������k�]l�-�i2*xq���q.�s�l�o.fYaA|�)��jS�),�k�LO���h����q���`_3��;d*~���K!��CZ�ll֐x���4Xm)�Xr��X�n�ZA_r��E�C�:�ƗϿ��m�����]�"�{�,C܆��_���锺�]�I83��A4H�����B��"�OI�O��7^�;K2x{���W�Bp��AA���d�g�(k������|�+�5<�c�L�12����o��I������!�ˡyƺ�Ըr�T��'�4��^�.F�6,�q������=�'���`�@�G���^�ӷ�D�OBjA�$;�2!Vr �#��P�1�n�v�Y/
&o�b;��uOG�ի��C���c.,LV�U����%��@YѫM\7ͅ�SP�?�0@�]{��5�Я����C�%��(�h��k2�2%���V[�3�|>IiOg!���B�=�2���[-���:�����B�L�3L�Y�����'NsM|y�8G,U������̇]_z.f�����K�4�"��w;�7o���	I/cU3(|��/�Ϡ�3����;Gn?�R�.��}�4fq2�B4B������e��u&�߸��	�K���Ѷ`�e�N����Ԛ�y��ǆ6�.�87M��9ۮn�0������g��d�W6�w�*%��v�I{�/�]��l�m�>�uc��'2�V�d�⃀Ah��)�m+�L����?����H�Ӣ=�N����*�gW��x75���5���,���E"m�\��hs�D~|9�~�k�ؖ]�H���n��x{1��LՙfDĔl���z6z ��ĕ�
�o�����9(��6_`2���eDx��x,KN��E�)x�N���"�īkA���W(Tg��YF�L�J_�	�ɨR8�J]-�#l���1Ʃ[/��i��4d�Y��"{�"��q�ݚ�� 1��Aҹ�S|&F��>�u�q��ν	B�Lݘ^��M��b��X?���{!�;
|$���B��?@D��^=z���^U�#����;r:��!������;3���}ye
����i������Y��60�o�$&$<��N����_k�P����@�d`ٱ��o�~n��mIa,���̩�񶁩�ڈ*ȥ>�D��ÿ@�"|��_��60�~��^��V���܊�|�WPB�����#�g�B^�  �&y����{E8��e5I�ʊ�w�!�5�^�����C��4Zcӕ�d/lM���8#�r���~QY�rP����G/n���zs��?�b�ʸ��>WO�
y[E�%j�#%֘�}'�b82��i(��,�yL8�k���h��ԧ�^�kR�B�K�Y�꘍�E�D���5��^ҳ�Qᧄ"Oe���S���1�
4v�_P	w*�̸����1��+��,��Y'��/��i@[�5�g`X��a�?S�n	1��	$�R1��GF��m�����Bq�w��8^���OE��-���[|� ��"�/�
&�;��=~W��+�E��s)k�gq��2�� h}�^�tWU��O��"��b��g|�E�G�U�0V���;�*�]-U�nP�'&��wM�@�#��m�*��Q��J���x���b��>.��AN��;\IHn��x�����ߒ�<v
9�Yj��șq���|�L��F���t�[����x#�K'ŕ�ݜ�����%�S�� ܑp>O��ȫ��Yd]�0�Mӊ�Ӳķ�C1~�!ukܸ+&_YLi��[��U��.���=���vX����ϩX�kX{�>����d�r`d�x����
���-vq��r�}��@D0&��9K�2�GW�/��rh"*X�@4��$����৷Y�Na`�4�R�,\25 Ƞ�
YRW��#�U�,�j��s;ۑ�����Zώ�@܀0�Z��b���0�m�:��OיI[�f��b��ƚ�&p���
�`����#at�7H�SGⅸ�Q���w���������zA�j<j�|�
)�cԇ>y�o �z���"���Oߑ�~]!�U��!�f<�%K�V���. ��M�>�>�� `���&���-��t��w& #���F®�P�w�{p}�>P~o�E�x�=��m@,����zx?]Q#%�1Ό5��6)G��D�t��
CŹBm����RwV�֎M��d� ��cBZA��4�e�!i6Z�>WmNp7��Ҥ/��)3�N]�n�7?h� 6d읽�|��P�vV�������	0�:{d.�� �TA��B:{������}Z�������o����O�he�ښ-B�N둨Wx4xψ�B�8?|� ���^8�*5�o�a�[u(6}��gd��AVH�iL�u�-��p�ꐳ����%ф�������#�1f�5�ee�GK�s�wɨP�}��?�g|!瓐�{���T�� `@����_q���%�v�-�%±p�k&���[����k�&��?zM�����ƀ_Jׂ>I�e��K��'ҺX7���Ŝ�/���e����/if�*�G�I���M��yff_
�|Ρ���s}�'�J�,�ӭ�b/�%H#����˄8�>JT�K�,A�^83ć2r�z�^'��Xh�����&�]hy	��(~�=�y~�:��B2Vs�Ͷ����ng�,QEU���>C�+6������rj�z6y����s�Њ'��b��$؆L!�/����2T� }ۿ���K�h��E���;�oݫ�|RG�ˮ3z�Zy/:Mcj�|�O�as����鬅$Fn�@4�Z��sQ}c��[Ln]M��RG�V�qd�k�#I�eI.�}�)����N���tΝO��C����������tTO�ܜ� ������E���O����k�ZM�N� �����ux�F�'�q/���/���ak��%���L�..I�(Np�Ĉ@@�0��(T��E���Q��_�7	�_̸���>�|�X�<�R�F��
��c��ێ��I�̦@	�&`��%���D�-$�����z�1B��gRHt�|^�o_����p;�iV�B�e{�=��AX;��<p8`}�sZR)�y�D[�~z=����6��6���mO����nG��Hcw�vR�N����$g��3a������%-��.�5/���U�����ZU�F�K�6b�d$Q=�@��Lhv��k$�yA~<�����&h������<�����Ѷ:� ko���'�������vkvL����T�eM2����<��B_!e50�(�]z����G�,9 �� %v��Q8����`>_�5A�����d?�Y��4�r�mq��L���|	>K�Ȉ���}�%~�ٻQ�4�FZ
ߑN�_=�X) (b���f	Ev�\���JO)Tc�"��%��^�G��+/b�1���A�U���,�Ã�>ꮇ�=��<��M(5�6�n�����$ǰ�mw�x
�E�Np��~�6K@���g)@����La���x��~�>�,�=��W|����D�U�Q�1�:]��	�H���D�A�X:�4�B'�w��n���+#��hJjt�Ҿf*�8���C��Ui�5�\�p()��.�8�-`�ֻ��5E�� �.��*��\sg_��g30Ƕ�{��	颸�tW��7΍�-���(���}����8�1O����n�����Ic�	5+ܑ�i3�����*����$�t��8�HdI������x�j�;�����E��+Ó�����h}a[�����I��-���R���I!���6Ax����:G��ܿ��yjʘ���L�%	��I����n��G(fF麚�j�j&����A1���4��Y[A��!�t������
�lctw6AA��@TW��3q����l�"�IO�GlqC�К�)㽛�A�_�(EX�Ҝ�7�O�&1q-G�_�S���1���#���m0n�|k���©�y����!��κ�S���׆.5��bn��6��̧��[1��9@�kE=�@wv��/X/U@�$�Ž ���l|��9��Ueԝ��4w+/�Gf�=�<�z�)A$��T�����|h[a��0������ui����~-V+F���7��8����;}�XR��HX�!���R�n�.{!:'Q��y�y+�S#�)���&ZX����,B�:�J[H�2&�Tz��;��{�5����*��C��r78���lI�yn*�{@K��N�0����ޔ�vލ���p�^����Mf�4���ͻU�=F��u�՟���e��/O��C���za�У>��P�ɼ �>F��}Yg*@���E��ǜB�}��ò�P��)J[�l�{���^�,t��l�
�� 4P+nMa`.���REW:7r' �>� .a�J
y���A���d�6�嬟4�:���f��J'a*|6 ��W�o�
E��i�����:�:ٽXXQ�>��<�9-s^.����[�h?!�'5������OQpfJ�W�����
A����ZZ������ؑr�;}ƅ^Mڊ�)b���PMwFߺ��O�m����s�B�^�Tsł�|)d=޶m�8<��;�����IOs�D-��r�i�'X��bW�ᑛ1V�(�.�8g�_1�S��M��H7	��X���?����}��z���e YR����l����
"����;�'�3/}:����]ό�^���>��).�5��@9����:��������.q��Z�|��:�ך��f�3 `�_ k���ݢ0���>yī�Ԩ�@�
��_��&�&mD�'��D�T2�V�v��Fs�+@�u��r���S�V��[�r���x_d[��/��;��Pd@�m*Φ^O�~_+X %��~���P��Č|�.�8���-;r4[IJh���k2�33*'������ţ������CP1�=�!F����9�]$��,F��S�~u{9܋Z�b�t.���="�Gm2�N<v�$�6�n�'�9y�8�.�c�ݠ�D����	��B��~����q�:RN��1,;�k���6�W�wC��ɔ8��ď�����݉���B
�	g|���2��6��]UH�w � 5 _B��U-ə#ӌ�J���,N5�k�:�l/F�X�D'�c��2Ct�,u��5�A�`M�/s����杵+xg��C�s���l��̮.Ly
TD3#��\�@%�oeVH�5�o�/t#�dr���0�v��%�r}:��а�0��F]t<�{����q`�O/ٸ�\��7~���2-z����hl��������W��QK	{||'��e܇OCj���?a3�Lg->``�|!u�F# 7�Ճ�q�������ޠ��|����}4n�m��ĵV�B+��g��%�H�FC�]�E�rO;���S�SRŶ]O�J�N�(�x,�QW��]V��q;��h�^�o: �Zz�])W�.��:�gw�[H��2=�P\R��t*�T�Ŀ2��V���>�0��'òH~��4��������[3E�$o�H^T�#B�c;77m�IXE��J��u�(#��zQj�l�\������&-�W�f��8�����UϜ���5@ug2��'���A�
Q�6D�Ȯk�M�.y��a�'�$(M%*��D���-D�e���%�`ں�q#�������[(����MtV�L���\4�L�bba�[�Zg�L� ����˾{U�A\(�
��9��J|�{���p�=I��#c5&����8��|!%�H5��n�k�]�_��܋IƈшG�S?У�>�b/7|*��B4�e��2[/�Ot��y�%ۃ������;�	���û�^JA���_,�:�����r^�lP~�����q0	��}=�8���s����q��0�a��(���}щkV��Fj�>���a'�7Ŵd�-}^��P!�J@�9���[���3�͂ʣ.@7���)���	���U�Ջ#�%O~��蕘�����%\dQ�`����y��]���G�{�Ǫ��&�Q͑���*��"_���,U��]��=��ɣWg�{�TW��~����s�*��)Y� $p���rF�
���o�!�l"R0���*Fm�f,��`cly���j����s�H�٠�mC�0g)y>k�}i��o��޹\#���'[�$[�˕��=ٵQ�5LXd2�s����JФ5])=�����f����.�X��ڵ�������>D�����)=�C�WE1�)��Sa�	q}[�C�_�nė������A���h
X��I�-�X%���b����(��7��h�{����h��ӊ�� ~�k���.��j=����ʍ���=�㮞��(�4x�.���N0E�zZzLL�j��W��jQ��A�����7M�d��I�&�F/*>��;B�'S���H:��᣿�� k����a7��R�3�瘠�zx�L#OEat%_ZT��/��\
�JZ��T���k�KT�h��Ƚr�M !� ]4?��v(��"K	 ���&ϊ���J|&����+^�|U/$��sL�u[qꥨ�R+n��TM�1�`�l�q��-��gD�c���p�?�6�<��b�(�ǻ�=�ٹdz�&Uxd�E�>T"�����br��?��Iq�.��O�J�#�Y���C��t���xR�-b�9� YG�bѱ�b?@�NMƹp�#��fW�,�Fw�j�8����5��\wI�X�	��q�I�:�c������]"�G���fg	��߻Z��塮k�D���w%��p/J?e�Yy�t��?r�)�ul��f;PO�v'W�$��9!���ó�@*�o�L�>�Fmح�+�Z�s�v���P��/]���<M�ks(W���LY�[�t#�T4��D<�mлl��r�t'3NR�ٸ�����lʔbI<ZVJ���!���w+�dɈd%,��"��¹�q ~�E,��dZ�'q�GMT�g�_��<�B>�^�t�����]�w���\)-p���~8��wG�G��J'�`���	-V/
5�a�D
���Ioz-�I�<��|�- ҪN��9�%�8���{�+m��ۓ~H�\�2����N���2S~p�:������?{*ŕZc��|�Fy�lQy��EFo
��xAjP�� �}�jK`;#��ac���AoY��R% �z�R��}��TW�lc��P9p1�xQ�>�������1�|��.+��� �u+��k����jaX��H��c��u7v��.M��{ލ��sL>*�Kʐ�ɸ�� �t�^8zJ7B/�P�$��o��Ώ�}�8ګ�tI�3Rv6��	ϰ����DX�IE;�a�����g�A�fl���1��&�PW��b��N_�$�q�9,f���R�L�1w���ͣ��g�6��ι1�ޒE���gwl���.�:,}1�� :�:p��1�Kb"�D�,�������x����] �֢I����U9qH�9�_u��@��+����[wc��$�pȕ�ő% =����4D������q�� �1��[5}��w{Ҕm�3Z���AAN�(֧��e�1,d���2|�R&<g�%0�Šö��Dñ����7����67��g[&�3 �h�AD#��<P��	��{=Mt)����Rߜ�wQ�O{�rb�,�U�㊦�� m�׏��.w�PE �>A��๫G�x�u6 s��t��b����{���C����t�;�/g�n�P��;�.��Y�7?��&|ʒ=�T0��mXI�d\��%l��|�����P�+*�֚�W�B���5l�)U��R<�8o��(y�%�*b��,>3�ls����;���5�2z�u��C�0n1��$YL���]�6FE˒!�'+��og�ƕ6qJ�ɦf��;���C�Wg���杂�>dg,��S0_}{���h@h�Ns]�����?�0���Gv
���)?��w/��Kk��V��/���� ih�f��ۖ� �<^�~�*��޽��h��R��4�=����Gʻ�b���V���m��X��>%��u �궉��#�h�n�.��
�.��X帔�ؒe���)��
�&U�ؓ�@�e�n��o�)�"�����Ύ�NZ��8KH<�Dq��f����e�Һ�'�*�s�_�؋ǎpG7咛ƈ�)�_͔$?>=[!��E����hj���U�E��K�?��%�W;�U�}-�d���5A�7�Ǵ��1atڲO��'L�l�@dN~�h�^(�Q���:�Y4�HF�*�^�=@+pM1������Sʪ	L�H_W.As�UQW#tqT��Y=�V�ɝ2ԝ�.E��)���ˌ�X�%�-[��UH�M�5��#�I ��{�	!���Ȝ�?R��o�h�"00��u�M�@q�4��[��eO{3l��-pN�����򨵟��"��t)C=�Ҹ]lZ2u�B���@�C�Y�)�]٩Fd��+��NEY����jS�����^��8nD]e z�Q�,�F#�+�`*u�D���{�B�Ͷǆw㢋샫�L����i!�S�;��Kq��QsА{ǆ�I�p"d+�O�=��>��w�����/RN����e�K��!��>J�@E���L7y�%妓,e]��_k���j��n�&����s�.�w*�A��� E�U�~�����ۼܻ=s�z���;��mi�\��Aui���c����Ω��3c��ҳ7e��1�����e�?E��=�"rH<b]��t��Ӆ�EzpLLU�~�<$'G��P��!H�sv��է�����uH��Hr
d-�0�O���K.�E���m�P?���G8NF�ٛs
!3[2�F�:�[YɊ�3wV�=Ұ+d�s����l�l�����~����>��^��B���pN��jXK�Y�OqF͛�ٟr��������v݁?�J�\�퓸p�qH�I[/l�B.t���Tq��v͋I�H:`�mC��fX�X}���:ڡ)H�u- u���}7��3�u私	_c���2^̍�.j�L�����(i+�1�� 3��b���e�ǵY;H�*���s-���E�\H���TR/d<�qwqM����$�lX<�ڐ�(��.��l��L"����&�h֊U�y�K$�uGކ(��6QRU&x��:"�Ҁ5�N�OO*�Z�lDY�1�ꝲ@�a~hB�4=U�'9WN(�$������%���?�|��%�b��]�ŁfZ��
�z��Y�7�� {Z��<~�K$o)����%�c�:�z�K��S�w�4bL��/H�Ӆ���KHџ���Н���RA`*��9~�x^|[wl]�3��wx�x�����s�
�����o��"C���,�@DI��6V��Ũ+�P-m#�J^��n�0�*\��,�)Q���JF���� �[���g�'*�<j���'�$+Qc�S��4"d��@�AS�Z�T���$"Dkw�Y���0�j7���n��<{����ν��{�;EI-���h?]F1����Q&	�Z��/�}]
��� ۥ��b��?�Y�=�����<�d�aZ�u\��<X[�1�*E_���hb̄hث=�� 7Ve���"@�a�8����~^�!�-IV*�C�)��%.�/�t�,PL[��r�S���1>��؈��p��֞��C���&�2�T���#KEYw� �M�߃Y^�·�L�(Rt̕�����
���;��K*Y�%��S',m�ւ�M���{��0ڰ�,I�z��-��^ >�ÿ��S����]i}���%�(�/UK�o����-OY��I������6���82���b�|����{�)��+�Jw�]�I؀��&g�tEc�@�}3�W܈H��z!�E��#Q�=�rVj�gY�ܜ��u��ؾ���9L�2�Y�{�i	x�^zm�U��採|4]2�3�9��������0��0��:�.+��`�~�EUa`���X�
�q߀Ld�ߌ׋�{#�G�n�4!x#�yy�[�Mm�#�uwRj�$�%�e#��0�M*s�/%�M����r�],��2��k��A"��-������9�.���6�E�Zb~W�2�
�Yǵ�
u�4R��o��1���A���C��N0���;��E'��wE�e��dK�֌�O��gh���8�����]Q��(4�����I�Nb'���B��b��L>TZ�
$R;��T}Zf�R��V������y��DK(�-��^;�>e`ȴ��ꗋ������k�:�ւ�>��)�
h����?�=<�`�FWU�7Mr�¡����bD�]J����dd�4�n��x�;Ʊ�mf��{����S�&��� �z����m�w\���M���/�UAډ�>0�_]�Mѧ�S��b{k*�����n ��O!���H�z���Xw+�Kf.������L�X�ojC�k��dO�^Ʊ� �X�a��M���Bђo�F ��=�Ɓ��}�}�&Q<W��!tzQ@�˟�����w\�n���n������jʎ��DD���?C��M|C;k���q`���e�9��^M���"6��2�N!���{̨R�n&w�jN4߼\�7�|��C�),�Q�B\�Rt�s�J���U����۩�!��}Ի�v�L����r�.��Oi��U�٥��j�6�mD��b���-=<�{T��KF�'��V>]�c�h΋�9f����So3��d)��sl�R��-��9�;{��)1��Di_�K%>�����}ްu����y�r�g5qI`�Cҩ�n+��5�j2��E��]�T�s��|�����L��̡pFH ����؈�� |.��Ϊ��I�'�Q9��C��`g��d��D���g"�M�a�`�]���{�C{f�_�1��5�j\>ZՐ �X���Ћ�F�c��x��G�i��n�����òfk��r��"fŋ���2*� �
���z�GOs=9:J?h@>R�G�}\��BK�>��L��������7�3/�@�CI�[&ܙӓx|�49��[.�B.����&|����3mA�f'��ڪ�{�>��Qj��~#,�#5��J�;�ݔ���������\\o| P���5̶�j����c�ai�Q�������`oėQ�9�����+# =(h���>�dx�A���~ns�iC6���iD;��`�����f�v&�[���/�� L=�]���޹"�2�BT��bC� �7� L
��A��l���ф���hm͕K�\h`�Tf�2g�˞;�Lc�'3��=��"�Su^�J�(<=$	�l�_~�u-z&)!��ػ���*�_	0�T(0&�-�ʗz㍫�
~��CЍ[�Nz"�D�ݕ9t�g#yz�� ��q6��)�i�`x'��-`^�%�a��EK�� ���6���d���׳ C�. F	�����0@�ń��ʺY�d���oC��;��O1��~���5Y�޺����+x��ׂ<��+�vQ�������~6n;v���ɉ��y�pڛ���L�Y�RDs�B���r�nP��$�S	��C����X��H>v�t"��S��z@=-�� ����K(���ku�'���aI�}��<�oL��So;���F��EE&$X=>!��:� ����e5�,�q���f��=')��G蠵2�M+|��0�qzD���'`�`Ht�ߙr��gTO�&_iɢf�.N�ع,��ZHB�U�ۀj5�C�2�)>�詴lj��-�"S�O;�r�5���`ʜ�q��Q�Z�*+ة�T��X�)�ty�ke��]HKG�'(��u���<K�n�X��%%�"�fE��*�j1$����h+�T��(X��/r�s/%s��}�����t�H�KM�.F��kĊ�~[P�ИOV2԰c�sR&��m��n���߿�b�R�Ф^�}2�������2����!\&�K�z�ծ����g��?9���J�˫[��R��OH��s^����\�iP�u�-Q�&��:F��H��WF�s��i!��Q��:f���k~�8�eُgb�(��{&�Z��D8֤��_l��0�l��:l�v��°OXu��F��Q�f�&>����x���a�=�ӬNpq�hI5
�F@�b_�����q�(aP?�$֋m����#4��]HK�qj�-̾��:����!7
���p&�|�Y
��
nE?�S.��	T��Tu�������Nsr�����\l\��n��83q�wN<���Q��&���+ɝ���+�J%�Y��!�*u�;���MIˤ���4=|v�5-Yi��DB͖��I�V�͍��W�?�$�#0��"K�����2�z�ZCnD��"ʴs���������'myH�־b.��}}���U@��oGz�M�!W�7 �v�ԑ��W}/8�8�m Q:�5+�׆`7�������-�u�K��Bk7Y��J����G3����'�.f�f����Q��%�z��P��xWBޚ��M˱��`w 0��	|C��D%XꝠ���Ź���������Gu���Y(<'�fM�u+��Vo�etR)-��������w]��V�<�6�eK�k�j\E�֬%~r}�7�t�"bO8#-_����K�]/��M�~kI~�*��7d����u<n<�R��y+��	%
�Vrs���A��!��*/�'�-�z,�QD��G����8���%Np�ίl�o�p��)Q̀:�xq�h��M�}�L�ʌӒt�9J�B�7�v�{� B�x�����)��ߦ��|�)\�G}j��7�6Sw��%��g0e�4XH������1O�$�5>.�.PE�{�]���8'F�dΉ�uD��a����e%�.�=>1�)kf� �V��
jnڼ�z~/�"���$iv�(��c��� O79� $��S�uxk�b��$b���ڜ>��T ����)�e�'$�VK���C�ED��20>7zQT�8C��[���nju��R�w4�]KY&k��p��_%��LU�ո ��*��Q�+�����H�b�s������9�P}^J%�HN��9>�w3+���
]�Ȣb5v?�]D�p�����к��Ak�jo�^���E5��J��f��tL�sT�М�I��B�nif�HQMm�>\���ytb���|4�F��]�UU�c�gmSS��c��I	�֙C^�G��#�z��`I�c������.�;Pαa���0�� �q�N|�-�Q\K�5�5�UG�>���r'��)%|�ƕ%�IH�*߄T�V@[�}Lu}��?
����XC��Mڊ�6�� ��z�E[�:%py�����2�-��g�ʁ��+থ&5>D�n��R���r6�݆�A&9�|���	�ǘWI���%IW$�c젥\"���#)������ޒq��{��h��3Ir��vdŐ��ّh�l��F9{M>p�!�P��&<���G����&�	�T�#Lk��g��m�%o]�� Ќ�n�iKمn�]�f�T��w�4�e,��i0����_�������cW���m�);��i/gF��nS4K��Vm6�-�F����wj�_w
0�hh���3��O��ʔ�D1&����]�Wb㧒�zp���l���,^�^=k�Dg'�� �٥�Xw��73sp��S_lI�?��0�v�
<YX�b��;�n���ƌ2��k$]��O	BM0�=l"���N]�|pÊ�%��b�]���\�!g�c�s�1���ȡ��E���+Q���u
ZSk��7���e�g���\8��@ibw�~��૨�c�x�b����p��"|Ue=PD6�ID�|Ik��%߉����]�[n�=Q�>)�*�C�1����>7�$"d/��Ef��a_D���OA]Z)�
X���mx(,5��։�d������$�+�l`D����6���g�	ܫ�5z}��� �U�����p�"5�l���tW{^��,��E�˥������Ao��X��5�{"����j��Bgo^�c;:��jyyKw}��y0	��t���bO�rf�(g�5h�M���H:&@��1��(ȀVZm�f�M�tX�I� U)�`|���w���9����Ga9�ri����dXM[�H�_{-V[Ѽ�h�~!���D�l��;����m���H�����	5�q,��Ҋ�+0�	�����yO�<�AKR���~Z��DZ�$9�̃��o~en������˸��+Y�1Z �m@��"����YҰ�[�� ��M��Qt����p+�ϞK�j�~�����P��h�F~-1@Y���7�z���,���*��|	vS��3�M�y��fT��+b���M��5��Nv�}a������q��v�������a�A<]�O�ɶ�2th�LѼ��"�ݘ�(R89��h��'��z��ȋ�E��>n�73��Cj9�u�Ⴇ��dV�?S�,���.��)T�|�)n�t?r�I'[��u8]ƽ 	2�F}���Y�^�޳R���ټ��fU�<x���H��o���Y@?i�	�<DhItxU� ���;�M׶\Hjj@ȎgʯW>���zII+C	�ih�I��ݳ���w��EYDk��3O�w�s)�0D)3P��w��@�9������zC��>x���J�p�g�6*�J�zo%��h�r�Sg6a<}��y}y�Q,2��-��t4�րv��$7�/3��/�}��GE��Y&G���S>�3!�i�|Pw���]��2%�N�}3�TK��By����uJ �4��/1�Ad��[iƉ�i¤0\�cz��I�<m?UT��C#n��a�I����]:���>���j������H�"�ݤ��!��G?��/�_�Jp��l�P��1F&r�Q�,��:�>ِ	��>���������}���@蠨]\�]��J���vǴ]���BuJә1��>~���m �wp1T=9ow��y��3��0�+��:�~�ǧc-�ESg��mwu���u�z���VM���/��쑗�K�6C��*�����%�Ρ��A�h����zwɶȸ�[�>t���S�x�+�I��a����T��*-�)?�?d�����	��tS4&Vs��zO�Tw˶�Nݪv�꧑����uo^�Zs���)��
�ep��N��S�� PK   ��V�<�ѵ n� /   images/b6c897d6-7294-4140-aae4-5fd8f682e5bc.pngtzT[O�h� �V
E��{�-Z���w�S��
w)��/��P\^�}���y�Y����ܑ���*��I�	  �d^ Ȑ?��ӳAj� ���������.��v� �B��7�:��$9�I		� �V:��<=��,��T���޷$�͑&�od��0#�G���=����Ok%��Ǜ6�6ǣ�푀����Q\�(���P#h,.�	BE�4!	\FJNVԩ�� �|8>;ֆ�|W��=~��"��@$�8?3��h$���ѱ�&�U���PF��ID�y�TOp��2�e�"�Rڏ�˒�b(�A=Í齐 ����nҦ �E>xK�Ә�П�31;	�xL�E�D�ø�7F)���ӲDC�{cG�U*<�P�W:ogW�����SW�̞�>�W@+�ZfC�i̐��ҵU>}Q��'?7����[��KA�Q���i�e��{1n%�� ��[qQ`2�
�'�:��(�^��{�Z>�!��;�SH�F��M���O����y�C���4��,D��ҥHU5����̹�)�Q�&m��KRr�E�1�Tu�Z[��1�s��>_�)9�D66i��g�����cy�B-��@f�y@�5�`�&�q��|T�qtEI�6�����g,ɷ�R�HUͥ0�:5��,��xKEL���벂ˑ:�"�.xh�P,�2N��	���4�����f E[� dkev3�p�x� d�F�J�ղ[�_0?='��vG�E�	Cy�ҩy.�0Ҿ�R�#���IX���-L�C�����o�õi��Q'�25�.�Ń�E�7�L���X{l�F�rj\W^���;^��zt�w�K��]�L���j�!Q%�kiǌ�-I�⊀�B���c	�p*O �(6ō�����6_r�j,2F\z��C��k�8{>����ї)��x91������{�(�gS)=�{��Am۳@��گz}���{X΄�l;�/!Ҕ ���ZC1C�N)m�r� n����I�@Qv���F�
�K�	^�_������P��H^��m?�i<M:~�|����������ĝlNI}�yc :1�"�ᑆc�Q��{!ၤ$P#����ʁ�Xkbi��p`:V�$��l�o8�<�#��'�%�'� 
{��O�F,O5&/��(��[�t)�|�1ݣ� ����0)6_�%#>��E����������НD�M�3�=�h�:���oE6!q2ϱbe'O����ؤH?*M������4��^��.������:�ajb�
Tꮆ1�a���|Y
��a�r7�q�S�'k$\�\�"�fڨ9a���#}��U��{J}�"H�L��D٥#�g��)]]n^R@Y {��U���"A�O]e�m�B�4<~�+���Þ���Qf
.7�&
�������F��|��gx����[�UK[I��dT��R���a�"w�X5�B�t�������� ��Ҧ��l���i�+���[)�C�C�C����X�o)��~�ߙ�)��W�*���V5|�CѾ`���ˤ_��yY`}�kYaE_����sN�?�Nx-l��fl&��(��ΚY�N�N�N��{+��ǔ���ήیNO}v�,y�U.�RXN��7����|q�]A�O�V���В��H����P�X�x�can��>�����7�o_���/��^�],�N�]���K5�k����B���v�wu�g�b��_7��.�:�pu����:��Í#���0�����C4�'��T�
c�E�¹��x�u��D���*Ĺ��mþ����Y�3�g��ϘT���VAQqU~�E�ȕ�u�5�:�7��˩��� ��_�Y6ph��2�2�5K7h��+s�J�T`��e3L2L�����5wiqّNrYƬԯ�Y˲ե���y�گ5����*���VK���,�7֞�9V��u�VH�'NxBZ.2T�T�qTK�xr^�x�E���Q�=.,n�>��ǔ["�Mc7�J��� D��Jb"�r�=Қ���d����3o���؆�����/Z�k�i�;�;B�R9j٥6!���;�8K������6��?�68c�Ǖ�&l	i����	�8�`>�=/�Hv,?vX�ɳ�ǒs�y�����;w-w�����C$�B����WM#�	�p����n�Ml!ʋ���A����`��%)7�$��Ph����E=K�
���'�v�9����W�}EOH7'/��$ǋ��A��n��u����q2yݻ_��җ'BJ����_�q]�q��L��ddWj�2KcP�Q�UVU+�K�]����`�����2�K�/���SI�����,,���8�ƞ�oƉ�wZI����2�0QA���ƮGb�^��rfPp�z٭�(�Cxە~2�0{�n��q��7�,>`7�T�g3���y��c7�K���� ���hԦ�/��_'���&i/�k�"c\��b�Y��+�/�f�v-�m��3C���4$�����ӓD�&���-��,`˹,}^���w�r�J�ͽ=�%��������vi�Bj��Q6!�����rS��kF�ˊѹ�6?+Lfٹ���_�>�<�d�`����/�Jcɤ��I �Z��swf�-��]�y��OMֳS��9�|lL��Ut�����/b^����>���O�P�Ѹ�Ự]�RwVG�����W�,�ѕw�������(��+'���U��l�����[�X���۾�g��o v��&�}�`�ޮu[���1�z:gxڬ��}ȷ�ZJ^����Pq����d喼0��������֝倀�|�3UzD��]�����I��pY}��ΜF�ު?ú�R�c�Zޘ�'_&�k�i�������Y��Ѥ�#�&�e�&_��A��uպq"w3�-u-��n>؊�>�m�}��!����}�>]Z��_Tz����k�`E����e�{�7!9M}M�>�/)�~(�/8���9lY�8&Z�kޡ^{;����A����t׆3g�BS/������t���)W�T�(���e�~ӯ���a���]?f�9���K������;��}�.��Rێj6�֖>4=}��X��i���v�H?�����*�|�)�,�P�4u�{���������5Q�O��j�W!@��6ߠ���ۉ$����������#п�߽�"+p����1P���]��pw� gI4ojbi*�T��=���b���?Uc�|�-��ѵA��`}�6�m�� ��ǋfʀYԣ��w�D����?� �\G�BE��P��h �?E�⿰�s ��02 a@��_�ϓ�o��%)��"�S�>"�g62�#����$5��Ԛ�.���V�n)^":0�t] ƿ
��+��?X��Z:n:*�B�����f�&��^�N�/�%��7w3�z��9�
y���=C��W7��)n��t:*�PiGs(;�F'�	�BE\�,�^������%Jg���$�����������b��)((�����b�3������؋�����E���������������������(ݿs�y������vrp��X���';��k���_�B��^�v�2��h�g1>>�����S��y��L��?���������a7��a׿������Q�2s�Kg1L���Ls!���)�eԴ����Hқ??�����%���. �@QFR��#`Y ��٬l��g������P���	�ېW�f�p=�����N:Mefs�T�>�g���0*2=:::��j���j���u�8�#��풣���p׍7Ӈ������y+r*�����5�KO���q�rW!q��_^c�Yq�?b}�,���d_���3��O��Ȟo:�<}����p]ǙJ$��,{j[�r��W���n�r}U��-������v�#�����C��1�GH���a�L㐝}�;Ǟi�
�]� "�]����o�*����|GN^�y�|�_�{�O`��WM��<�a_%��֗�AW�\67J~S���E�E	�񼫻q�ۡO�F ||s<�4��4�|�_�΢���Z�9'�=p1��J�
4e)�J�K^���e�E���\�o���)�ҥ��jSx��`AN(́B�mRM`��n��#iC��vg����@NC셒����C�}�]˱�����x��Gm����jv�_�ݢ�s=�ӯR�ظ�N�;����.4-���	����߉�J�VZ}�V�����{�4�폷J�'k!a���U�3��v4�����jiR��Me���_,l��>��1ʏit�sQ����Z�W#�W���v�iJc�H3%�A�= ����n�*���Q��N=˥��AV��0,:��"Q��K)��1-���J	���<�?L�6]A�x]Ģ���lpM��p)�G`S��%��;Qx/���+R_��O��\��ҵ�&�ߘ�$���?��D�S����ؒ�B|S����tUrhP�Ȑ~� ���!�-��=�ctx�Ir/e*��1����Q�er�LM|�~M��S]w���%έJ���9�ׯ_O�>^6t����r�;�W��b�=����fɚ��_y�J��R��[�b��6�i��&�2����k���O{�?���O���*�%��}����]�lp#M��p�o�M�l�������5���+o�=��F���?���k6�8���w?�[N[c�h�)��8�|G�ȓ�K�I�{�Y�f�Y�7{-ۼۼ�}�u�b\E&w|
��^^JRm}���w"����n}W���/=���j
��`�T��Lm#���.�{�.UB����~�~�	<??����5f{8y�E�H3�'i*+�#��߯h�����i�]z���l��k�?�5�R[:�1[���P�zr����*��ha�)�d�Gӧٛ���C����Ԗw����٪J"��Q[�F�7����_�WM��,�+3W{�.F�m͊�E��ć�������R�Y������:$�r�ɫ/��Vs��Ҫ��f��b� 3~�ܠ�G��DS�l&�8�ܝ�F�~9�J�Y�y�!W.K��o�4hcϵ��.=���:�	�++a�|�sS}�/~��Q;���k�m�X���+��X1<��+�V��|�1#�6�Q@l0���c�e3�Y�%�/��-���+��6�(�_��O�G��Ά������ϲQ,�fۙʽc��޹W��rV��
��p�͛<}��ͩ?��Pz�p}Y^q�G���ep�~����{�Y(�r롩�1!'Ơū-�ч����X�I��H햍_��->��`^u=�tR;�3�(��2K;t�k����W�Uͷ����ۍ�˝o%����}�d���=��'b\s�#�?.|?�ٹ�qP�5�������x�W�NJ�$����V�Κh�I��A8�k�v�rѺ��c�p}�؏ƺ�Zyuue���.֌��g3o�:5X{�h)*� �8�P_s$�h��wR6�aG���	B�TK��Q�U�΁�M��#ydM�4��5.�>�e,�h�Pi���N�a����j�m��v���GC����ܷ� n�����*B��w��z�;y�:g|v�������r�6'���K�q��O���I�<�m����݌�����Ъ$mM#O���੧%|�l���jn����4���M֣E��P�pڸc^����Ŷ��ļ|�.\���4��M�C���A!�2��T�~�Za|0��ԕ��$Ʒ��R#N���(VB�<Q�$��H������p�C��8�h���z��݁���e�w����V�L�I�f�/�I�Q�ƛ���J���enti�r�"&~*�kQ�L��D�|�7z|�/��p�G#���9cO q��㍉��=��ZW෡�=����ٓ�s�9/��Ũ�|f�΍r��?�K�O �Qڅhx�cM����0�V��i���޵������Dq����1��62�]��(��X�aS�G2~�?6(�k6?~I�T ���	�h��{���y��W/`����!�n����×~2�з4�'��sM)y�H��"}�T3�>��Foh� ՞�W{%��;m)>�.�
�|ڱ�دݏAvժ�b��DaVFzc��*�$���ɶbe�[��C�4�#�`�v��E��~=؋�B�V;����G�p���t لFE	�(F�a��g��xС��������ƈ��f�BN.ያ Q��x9�ϱY��L��ZDƠ��v��,���b�y���:�d�s]�����	�-���*�0z�
���\��#���j ����a��U� $���I�"�Ư���Q��p�&���2&~
a�K�.s�_�mIQ��=�:����y��L�S:��}b�[���%�g ��׍k��r��� /�/��*Ru'>��4 ���UN���TK@?�s&P|������
�-,,^��)
	
֭�
����mSu���@�k�W3���v�*e>��	�`��h��xCu��K#�ę�{����)�7%��ٗ�Fb�� ���ә_?B��������c��
ns�ӕ	�	�m\�6W�ۙ�ɭvbC%xЛpt-�Tu��8@q�F�9�#�������}��fo��q��ɟ7g���<�]��Dn>"DP�X�,U�
 �,�#�/F�������'6��.>������M��(�`�s��X�%�)0�8��i���Я̿�j�9J<nϏ˝�%�a.�����������3�Us;&2Z��1��폷��b^���k��e&
�K����GHE�Y� ��Q��{�e7#p�j3�v�+!h9&�N�}�?f���+7� m*�{P���
᷏��W���4p��hO�+k��o��YB�����Q	��,--b�c� N}G��L��@f>Mfmr0�>�oM� �tZU��߁�r0:�\5�&�����K��A�l�:/m41`�\���}~�PuRbk8F����,���x���}&$ohr�Q���&���&=��t���4w�|-�$��O8�ڏ'�����������I�n&w�2(|�+�2BYXP��A�dp�/�z����m}���[���T��D�p�)����|��q�ڟ�ѩ�d�/�J��1Т%E�D����G���N�IM��Y]�,�F�[%����lt�F�RK�c����@��YIT@�ɟ]�.��n=�����KH~���5
��x6�����!�&Bl#�_nx��+º�U��<����b	���q-l#ER��<A�$��y��{��[T��tP�䚱��r�������v��~�������x!YѨB�X��+�g�f��9�]֛��e�7���pB0=+\Z�ɹcE������Ƞ�l��Bje��>PE#V�i����"rf`�%m�8�4����y�' ް��d�-�.����Q����&�s���"@,�2B[$%��(�h\����0˝�Z�����e��`9,zVJ��y�[�7��%m� XJ���&�v��̰0�U���/]�q
��C��%��^�|�s��j"Ŷ���b|y�o�#2g+��Tб�YD�"W�R�	�����m�H�c��b}x�#����p���|�l�o�ã�x���$lU���vlP\+��tY�r:��x:p/�;;u�N"|����U�N��(��)ͩ�����ς2X�=ɁA:Ϸ��$�t���!�wR��\j.�O�
"q*�ӡZ�آ?�P����'zC��J&��O��f|��RR��*pmĊ<Kl%Į��P�q�ㅎm�z|?�
�MJ��z��xa��h�=?� ���Vj�c��jj[Z�������?����G�.TM�\]�0_1G!�ig_�P�D `f@mw�4
y���z�N��ul����K2Ȑӏ�K���Ӽ��_&.�w�wGQ.��9?�@3�D%hZC�h��7Q�,+`h���V�n�x� �Vه�o~AO����8���~+!��w�I���A�gVl�=�|�3�<���)I|a̖���¹�����0W���y,$"!ݙ��K��7��\g�S�x] $u1��nZ<�͍������xRY6n�*m�X���̺�\_�j!�9�y ���^���'����v��
+��|�pWK���-��5I�kI��;���$� H�]�C�;/V�-����7m`�)���`ŭ�({qSo� V���r	����X�K󜶠qQW]v0��'���-sԞ[Q-�O�9l��5���$�y�A�\XxD�}�/� %�mn~v����i�?|鄘�t&Z�8�� L�#D�|{�P���["i�;�;���_�,�K��lO� �:T�n/��jt�jd�TdC��"׿o�Z������ʫ�g�DE!˳t��Ŝ������#��}g8���^��9/�e����/@�Fx�Xv��9j�T��kswm���F�'���˾�$�K|v�~t�#rei�j�5����&«pu/xA~���Ϣ��	�w�OyM�%)|�b�:��'p-����������/g����̖��xX���g8B����b����L~�CY]���#�,`��-�n?���6r$���]�""���D�(��sN�y'v��]K`�G<0��c-Gj�	ܞ}�$B�0��)��P����IH����P�܉8��eJ��� ���O����p�G�]�ۏ����/H*)jU� �A�I��fNa`�4�$/R��;�m�����~@��A`Bj�S�e|_�1a$�ΒTw����:Z���#�����r+�Y#�n��������reC�rQ��?�`Y� �vn�������m�?-e��v���׺��eR��J�|#����뉾D��G�i!�;�2��T�b�������8\��D3�"��d���������6T��߳�]!b���FC����/_,�,�Ph��_J<����E�+���gby~��'$3!BjJsL������~nv�5�!ʹƪ=S�Y�#Y���O@߫��ɪbbҤ�]2�fe����Jn�7�7}?8���}f��VY7Wx���f2oE���*u7�ȴ�%O�L�s<�i+J,�W���O�H$=�S��c(�_�:frD�|5���O:��0`/?__�:�KMk1;{룓6�])*b��K|����-(�����f\�ɀ���S&G4����2�[�@a��x����3�Io�S��[�%� ���&��.A!�8?��zȓ�X6u��"��s����p��c��as��Lh7o1\9t�Ǐ�x��ͶOA�u�҈���]��V�;7�$�f��(z���|j=ݷ��h�tjk$�������5k%�$���D�a7=Eq�;�2Ycþ���'��]+fuF$�p6�ʻ�@�Ixа֛e��+�/?H�yd/��cgG��YBR)_��U{tx���Sδ�`Ď�U ���2�Ag\�����S�lH�������%���vu��b1!V?���՞�3\��C`f��9���y�U�8���.GX՝NQ
�&��կ���
q��\Έ;`J3�Κh����r1.��V���2NҎ�L@�
J]�T61�i�Q-MjO�	�LdH���#�Yd2a�d�-�sTK_�inZ��.`�=T�k�gc�+����1U
�~�5md��I��d�(���$����DM�İTw�Z��:!��q�jMʹ�`��L�p��7���)�43��G�.)�{p���������[���!�rr�N8�W��gz^ zW�����Υkc�����9w�zL����Ť@���ŪW�C˕|�|.U��A��رn�.��U����hşa��[m|�6G�(*���џ���2E_-����H�s�D_ϧ~��N=���.�ɮ�W}�c���*����-"�cԞ$����b�s�uxq�a'�����#�LC����bE� Ԫ��}����?V�s � ��YH 6�¯�H��*ܽ��yg(G�oU�'H_�+p�,Ȧ35��D��&qT��g�4����%-�����2��I?�~s���i[�j�C1(�c<��0���Po�ܩ��.J������[s��8w%j�$u����=���x��g����"�@����RRb˷4�!-��G�#��n���-��0!��Hw�E�ڢo��6�R~����^5n2�Ժ�/��eY�w��-�?�6�@��Y��4Nn��i�)���RU�� 4\K���4 �v����T��5��d��V6H���*��w��::CQR��6�kdc\�7�\���%�{N�r\ȹ�G��w���8�������.Rb@x���<#���&r �@3qb�v"b��~����9�Ɨ#���_ha1�+y���F?ھ�r��+i���b�Q-��������b?����y�`���QWsǪ�c5	t6n��hV�?wP�%�d�dCM��-1\�h��S�j;F�O:4F���pr7~�|�w������ƍ�(�mu�f�x3O��랈a��x<H�P�|i#Wȸ![ksUf�n�����z-1��<��B�6���z�Ta��l\������J B-��F_I��f`��k+��}#S}؝j��?_o[�e�iȐ�Q��O��xbٴ�S=����K9r9ÐS�_	->�e�\��!_���6�)���a|}� �_�֦�ݥ�dG��=���E�0�]�s�g���m���M:�����0E���/��x��@u*-���'r���Ƣ����E�p7<D����g���c���@��'M�;�\���3��I�����Al�_ֆgxjh5������W��\��x%q��G�Q~)X�p��J�Z2�yR.|)��j��H�� ����K��(p���Y�+>"v�NA�w��������e� )g�p�Y4W���Z@����liHv����Xafƻ�d�)
ci�c�/�Љ��#dqr{��WG?��=����y+�F���Вzdv�<�C�7��U �p}��A��o�=[a(5!�|A~b����+
�{z��$���|��T4��q��K1ut�8-�p&�;�(���ѭe�1{�ds8S�H�4䷻rGU'!�g���(.����C��_[bU�z�e��Kj��gA�4<x�T��2MW�X�Y�eDL�C�Dp|��'�+�R��1WXC#݄8�n �O��T1Q�0	@Z
1���%��U- �z ��n��?���3oB�$�3�&�r� wd��j*��%��T�`��<g�R�yPx�%",�
���+M�����y��)][�-�[�}>D4rĶv�)C�:f�V���8����%�9���������!DH�$��Dڮ�Ţc��p�*~,�9x��-ţ�Z�� ��I��f����Ǜ�*�׹���#8����" �y�uIV��-h��	�W����[�=�*��Tڰ\�I�NV��� o[}�P��P�Ou����у0p��?#�V�橓�+���#�Rko��|V_�~�1n劽^��
v֤�B�(.Hp���ϸ,u�6f��8yK͘x�c�n�<�P�ν�x�y��O���P4�-�PWp�ڈ;'�'��oWG����}�0D��������;��fa���a�%��Q#\��d�u�,SA��^D�I���kI��0D �5���Z�y�u3�z�`c�F�*����X�<�� -iX���`�9�T�L�
�఩K>��@�T��R�@����A��؏ �E���T����m�P��Tw�29G��c5��H�K�*��33��"`#�KcZ��Iur?�A��_�qz�>>�&��o� A���������n'�o�T��v& QFE/CY#:��֞HS*$m�Ɛ�L�I�C�z+g-���֜y�fls+��J��d� FŶ��*���"�j	��m�<�:�*8.Of��8�C�'�ɝ�̐�nKw�� ���q�:؏�'��;�q~����Q�"�m搽��U���GZ��$(�EN��@OV���x������HI���*8���y�
�c��%�g�U�QV���V{�sz��`κ��Cy��=����]��Jv�#s�	��k�!{���s�i���R���T8�u@(2�-�@T,d{k��Vl�+��|ҏ_U�_7/�ߟ���$Lccc���fZ6G�<b����[2����S+�ѻ-*��(l�f����=D�(|+N����C�u rl��>�{b�.��N�����7A�m̵���-F�_�^^&��$c�������g���Ԛ����+��G)b��V)��LW}��0w9�-�*�Q����{�?k�9�}���4ii����s��)��0�ޣ������&�>F�Sx�"p�e_�Jm(s�s���X������}b!���_��J�p���Sy��6_Uإ]�h��0���.%��e�3u���u�Es�5	�f���%C�xeS/Ԧ��ϴ	�l5��X�os��Z��m��0�xY/be;�O��m���ʥ��� ���U�;���;�gӪD,Ӏ� .�$E��eF��t�b�-� Y���3/l9�i"�o�>j�����p5�O'�t�X<���N���8Y:�����������w7]�}�z42ɘ��e�p���ux5��xp�\������7m
%��3�O�Q5�wbᬶ 3]�a,k9��pnE?)�U��������H$��u߿%�W}B��1��L�͐ÄtN��䡴ȣ��wK����d��zZ&���Q��j9c���Ghl��`c<�xn�¸�jHV�&��v��j��S*��y=�C$����|d���ޣ������!?��[Q�a>vT_S
���A�Ϩ8�c�ֿRnm_ʐ}1o��M�6ae���`⭤+����H*�)Ys�=\�g�v�X��cσ��>G�%�Mq˫!;�-��E���W-��:k9@G��V24����Pup��}�L�b���w*�c�ab(��&qM�Qo%1���O���L繵F�
�>o!�&�e��ӷ�vX�A�1؉3�ڕDE����˩�?M���Щ��G��!#|U�΄��h$�udT�Tei��%L
c��p��6Ztf�%����
_"�F����]�������OG���h���+�?C�(�� :.�0�*v)��|��.�P�R����@�����r��N38�	�j�S��G��,mm��yf,���9n�iS��%XP�7��'��t=���DQ��//$?cG�K��4�
��]�L��y��m��[�{����2w� `Í�Ѭ������ a V��#���J 6j7X���̮�"t�d��G�U�����������o��S�K����s���E�P�s���W/������&ƛR���!H�JH�P8�EpP�N�:-��m�c�|Hv��I$�E���R��_am�*��LD����8ݯceCh5#i��$2�?�aU�^ϴU4�����1��ىW���A��,���p_����!A�l	xP1�9�\U�����?��8�v��2�(.Uڅ�wP���?��,�z�u^=j��!��6x���.ۥ��(��{���-I�1C
0>�/�sL`���.�<9{UE����φK� �o�0#�G�^��3����6A!�8��V�rq�J�S�Y�t�`�s]<��M�|wIH��3�u��\Yr����?�CS��hվ�?O��+���?G/�fロ���k��(��9�5�LVk���3R��K���dH+�__��Ϣ�Bj<�73���H�F���'@�Q�&֊o����ߨ�WX�q�Flp���D�z"�R\'!A;�'8����b(�W;w*$��$D!�j0������s��ֺ:b,,��b�<��WW������F��X_D��"D"��xq�8����m�3]�;:�F�~m�gH��o�d�:B��9��� 	�p����[�*��kr�}���o����h��3��W)�߳�'��(dҊ�Q�^Px�V�O�!x%H�S#���m�4�
�T&���O�y_@�f�:��@�<��%�mZ��fJ
z�>!�}�E|���j5��2i���4�׉L_��'6��g�Qx�7����o|��?6��)M-	���g,[��
 �%�?	���oD�
���m���2�:1����RFy}R*6���,A����~F�൘kL�^g#�l��D�t�v�p<���%v��Z����׍$���b���eV�pH�q��	7� ���5�MN#�ݗ�9���� xH֬b\Ua'��d0��&�&�u;r9��?�lLE0��Q�l  b�/�D�}�7|�^2�
Q �ٗ?3GM8'�M�D*�`�Z񫮙U�u��*�Tߠ�?9�r,nee&��͛����*�+]+�G��_���F'�տ���t����)W������ka͜��q�>�[��jI2��k��@�v ��ihT�?��z�-/�&�0L�YN��p8�;Q}��>².�w�����ik�}����`�(�Z������'KS�8K�x��uw-�g����Y�72k�-��֌�|)wBL�%�N!���އ��������͵k�X�N/Tl��.��$Z�b��i
�Q÷���u��z�ؑ2�K8ʀ���7�����6��΃��������A�8 Ԝ�D�%<�w�4֘�Mo�;V���C`Z]�<\�o���%�ζ�/��_�(�4]���6��=q>��l-�8���t�f0 Ⰱ/�L�M�y�QU�����,*��`s�I�P����0�sd���mR����y+g��J�`��/�KSo�s$`bŜ��|B��SQn���	|�k����y︼D��'2nt
���T�2.X��~�\m�7�&�����n�B���DBrY�P�^P��(6��+UY���ʧT��J.�jK�d(��m�.#$�0��$�gd����B�ՕR�#��ÐRN�W�lK�%H�t���2���pu%�$U-S����DỞ�eԗY��#)԰
hm�Q�ׯƻ����NP�o� ��⃼Z[���[n���-	2���Z�I|��BAl�ho)�8^��� ���P͓P��+6i0�&0hV,�?}J�X)"�	
��۽<Z�>D'�N|6�p^�U7����j*��J��`��C�E,�7!�G?
)���G�A�Ҍ�dV��e�n�ԫ���(�,}�d؇�`#7�����pM�7�^�<�ax�Z�2k E.���A�}�k$������X2�2":Jd>X�g�n8��O��@��^V�^`��4�d��N�,c�|rظ_�ݔK�i	�w7m����X�M*M1���r%C�e���Us'
�fy����S��~p9�����q#���=�ۣ;�?FJ���K����Bp��u�X��#�y��ͽ��Î݂�g(&��K�����N�W7ˁܲ���	����8wtM<�#�_�������t~^Kj|@�ߊ��H���L�����I���#���A�����NI6��z�)�y����T�Q�t�;�R+�P��$C5�,L?!ł*=�d?�A ]�\�����"�r�+NFlR/2W��t�����H8�qSW�;��+���@�*��^�����H��1H^��̎T��kv#���"Ǧ�"� �Q�b:���	�����3"ll��o���\������h/F���K�˂�~�	�-f��ic�_+���E,I�����/%8�T����c&؎��L�+��a�����N��%7��������u�Ҭ.�d���_>��-����~A���,x-��I��K����wrp�b&B�Y!(͵�v�aP�ln6� ť�����s�����!��ldk��k���49c���{(䊶T�P����yBS֒	�
��"k(�v����� ���v	���'R�&����?���W�x�y��I�����n`H��X���tI�wD�"*TNJ>t.�iP[!�9�۴h��t���R����ܛ�n`�>�%Q (�Z�5Y�Y����+e��Q���8�G�CM���F��fK�^�t�H =s�V��<��N*&�Q�D���"l�1�h�㕜��J�#� �	��m�b��Xl�$ �H'�������a��Ι�y�Qߩ�E�~O�g�Xb#a��w5͊	;h�7� �$��~4��*�I�0�>��q�h&��Yh���Չ���$ݵTg 6`7#�Y��B�i=�tws_c>Hf��P���+�-@����9x�c�s&���.%c�@�"��!�䏤����6Ɓ��!�@���]��H;6-B"�S �)R���7b�`�����!>�%�iZ.���x�QM-��@=���3��Ix%�]'��Q�".����u��+�HɌ�)���-	+���op���M&�T'�:�<q�LvM�m۶m۶��n��u�>�w����w������^!���n �ț���b��O�PY�VvP`��oH��x� ��*���Q!I�a��"�qvU�X�!��.),˙�����Y�E7(o��'���iG��(X���o]5U�?�cu�.Cs�	�=j���163rN���:��LF�`�	�:C����q�lZ�%؏�&�z��8��A0s�lV-��B���'8�ߑ}�������^d���b�͂�яao&o�!cD�h�A�o�����?:��燅!�n�
4�{�Ҋ,/7ov+GfQ��f)�3(�7�q7?#�kK�A�_<߫��<`�y�YDv���.|�>~v���1ʫ� }!���[��9�y��G��v��v���3�! ��)�Ή�V���GNP�6�k�� 
y�B����ҕ����e�f'X�z&*ĺ�@�n�b���cC9������F\��K��@������6!Y:,��R��$Z=�?��XǱ����A�" x��9�O�o>�
Q�� `>��;J��q)�{>�&���1f`�����t��*��(��kH<�i2>K�e������)�;��Gܒ����f��.���L�fYkj�1UJ,��w=�*�~�v'no["#vP=�%}H�fX:u�w����]�	�)��e�9+A�_?K�SI>�H p �� ����Q�T}d�$1DLL8J,����$�҄� 8&.GC�WZ��_K'IBX�4"}�[�kFŤ?����"�2}����y�HD�c��p�1�C��
��'�uX�w��F"lM�����^?غ�34����$9�q��Q}�2�E�M!�tǤ��c���Nұ���i�*O,ϊC�;@��٪
r}���!��Y���� �dt�v ]�(T�ֆ���9s�_s:|��{(x B���c2e�*O�{��l��%�L��PN������M�)��+&�A�������������ϙ!�ɶ�����"���'\W5M�4����}4��)�a�JBDz�f��b�6-XV\.y,B��FMp�L��8�6I�(��Jݺ7^o�f�l"&�,DY:�'�,����E꣱�+)�tGU���[h_R�~�q�=aI�.]K�{��Y���b��W]�`芔<�������=+꯯�݊q��|��W��'�F���]�*<�B	�g�t�=2����Ϥ+�}r��P�n7we�>q�k >��#]��X6�ۂyP^��0�#�菄�����m�E�o�7��d`��$�B�a���
�yrlWˤfGGj�2+�iB3�Ȣ��	��d�f�&��r��
�����<�r(�Ľ��$�̀�GxQ����6��������#�b��5\�
9�(C��!o�q�s�<�����Q�d�>E�	��Q��̨0,�  $֝d'ЊM�+	�g�L���k�#�
�Q�Y|y{���w	���/֑!��$�d����,���|��-81|q��0�x�	#K�w�{�ƻ���FԓP��F���C>�s�5��c]G�x�Оb	�7���k�i �B�a�a�`H���)~^��_�6$�#t��ܘ}V��3$�&��PI����"����c;�Y+��Qi��sGKb]φ+���-B1�`@���!Kd��B�;,")Y��o@a^���ɘ����=��^CC����&���?P��i�6�N	��l��s� ����_���IU�B�E���ڤ ��R�� �c\�_!T"�G��>$�@m�O��R�@����u���Z��p��!��6� řBca62HB�%����%��q�3�,����n�ڍ��J.�G��9`��/�xɁ�k�5��(��	6�6�Y�b�ʓ�!^#5RT�з�H��R�L:!�
�}�fkß����aP
q����8��%�yG�[%����G9���Xoi�Ɗ�#��BK��'���_un�K-0�`��G9�E@^چK<|9��K�D�p�v���c�����4������Lom��:�wQ�D'ē�W��Sf� �YE�Q/��)���gmv(+|���� C�.�� �m��oϠ�)sӞF,2lH�Ї��BN��/��$aH�wx,��PR�v`T���+�d�g�.��v�=gp
� 9�o�6�$J6�(����~�.l$7����O�m�혬/�b�,̱��r�L���?5Vx��"�J8�=�8I�ExG�}�*��T�������}�@e�#ל>up�q]�Ah�{1�M����-����m��I�>���Vq�ZD}�EuZY:*�Y�m
+dd\�����/�����_�O���+Fm$#�q?������q���fT�_#gKy�t:�����(}-�Ы��E�QB�R +���އ$d������r�PRBV�T��㐐��O�;�;�ry�(����093��oFFtg�(=$�d��=tt6�䧶�5U����8vwj���p�aE�'�u�uXtx����-�QI)����9�;2X�
��>T'��.�e��5Մ# c�K�	�s���U4�#M�ȱ;L��\sN�B_��#Χ�}�#����.gA	��e��.NW�
�<�}Ń�h��D��;zV��ʪY��d�����?��?�M��}d�N5
�����K�f�%dt!#-�����<���$ȹt3Y���)�>%�7��pR�d�`]z�U��f@��{M�h����|��pu��眛�Q�� �wQ����)�~�mxc�r^)�e����uh2����� 4��*��:nE�iR?(*	&�<\� E��h	8u��f� �`�8ܪ���v���O4�ڡ�c�q��Ӫ�z�Ip��3�
3��i����]͸�8w�/���5CQ�]�����`|��Rv̤�f���q�":á+w!V1�����C��q�I�Q�\^�	7=o=��.!R�9>��Dd�2Ȱ�PgR���$�P�~h��/�Zə���pdq�	��h!p��F8\Q���(Y\氿	�{̕b���*�e5�6��a���O�����G˒�7�or�nɸ��M<�e�i[��!J@A^RΪ��~x�h���7�y�%n�.���t��D���~ڐ>1֪�5Oe�w���z��zw��.��+���,2u�X���a9��'��1n�ɺ�7�L������n2�W�F�����>l!ۜ��ټ�w@��?4�VN��`��O$G����L0��R�}�j>T��!d�.)	��j�-5��j" ���!�a�F�!^�R�2�!^�gx�@
�[:,W4j=�)�.2u]^^njiI��j��X~㼻���E��c6}�a�&R��|n+�Iۧ�t�6���+"�3�I���1�
�	E	���H!�CR�ú��(�v,^�72�oC�g�˶�M7��\��S?φ�og���s�7�v$����~���Dr(����a�s?�C��C���$�0�CJ�U�o�\u�e���Ľ0pl~�����'�ɺے�f�4���w䑍�
s� �1؃�h~Z���%�B�2zİw���PXм�&X0S�qպ�Ƙ1/R�.Â{��o̧��K�{v��������fm��H�5�k�m86�Ɠ�% �K�=rT�/����:WX�ѷl�j�j�s�tQ!�p"�ʫw��&�ގTeL�(�>�~_���a)����/��kH��2���Il��$����%g��I?=�=E��=�*�40�3���4���8ĺ�K�ݥ�Cqxʸ$����nO�$��R��0�ڳ�J��)k��&�p��r�g�(���?W��&�|�����@ܾ��5����ܻO=��8P���9}������|�����`���j������������X{��v�j5o�8�����9�A������2�Z�[^�?FbY����Ì��m�}o�2wl|)�锻��~��=���~t��	*����)�o��laFM���C]�vk`X��uk{��Q˘�t&/6j���S��S44G��£@���ō���h6�b��"_ə��waO�Yo��%�O���^��w��p�!ɘ��]�ћO�"Sb�!A!�K�CfC�,���)��n 	��a�u�P-�I�*XO!�$Zǵ���Æ�>��w�/��EMv�ւl��k�rF�׹�ca�S���ه��Q��K���[������u_�w���1�^ܪP�m��tM��k���}��-�G��0c��8��P��
CϿBje�h�&��7n_�����r�;�$*��{�tP�{}ϛ���cx7ޤ�o�]V桌�_΁>\��;  ���J��3��-���=l��X �c���Ӵ�q���ń
꿵�a]&9��E���w.�ܶ�f�` �[��{�Yo���rR%:b|����eXeI)�-|����!:�@���bP{C���V�� �^s׾��^|��<�T�6@ݻZ�m�q�� �W���ٷ�)�io�k'���� }�&It��I���#���_⪴�\�Sh���\H[�u�����Q%�rTōau��j{��_	�y���X�6W紽ܑxbS��� W�-����&L�|���eCym��D&]&���o̽O�\;{��>���_�I0y�M�~�a��-��U�څ&7�
BA�.ܑs�X���^�S��W����%�"Z	=��uL�kn���˻F�X����~�>������v�*x�v��������s��6�{-�oJ�&�Y'��w /��ϴ�x��v}�yB|r�U�)rv�u1����q�xX`ۺ��dC�F���Q=���BS�
�ai����Z���4�!W�����a0����D!f��X���}K~�3��P�� ��n�B1ܫ`֎���%�fw��+Zp��h\�a$�-��,��qV�ǈi�f&����Xf��I@O��=���v�#p����:QK(uX�l��eu멚z]T6��F(��}4=uJ�b�#�6\�bv��iś���qߖ�Ή������;������fg]s��"*�y�.�#��z�xLr�,�Ʉ�g��^w�B7t�N�U�΂�?(���ly�Z���d����6k"����ʼ�t�v)[X�l1m�N����RO�A�r^4��������tT��v��/Z�0s�?�������Z�fW�*m�1�������ϭ݌��^V&ŉ��S��Fi�Fz[�:.�u3�#�[��>�3�� 6�P�񮋶����×��A�I���W]��@n�uv��J\��=��x�/�>k}@#P��/t��m�b&5f򢃵�E�m�{wY�3�?杦���H�`��{�g?�A~� q���q??���mC�L��0>]\���\�˛}m�BKH�^'�]n�}%��C���	W-��}D��F��F�]b�kJ!��������65I$R �3"�l*)�C�&%����I_��vA�=�E��5a7� ��/k�c���Qe�RS��X����ق��h�{V�Hk�/�p39������eEv9������hY�m��׫Ԩ�;�o��d�3��Cc���3��t�Ɔ���'a�Oۮ�������0=\Q��K<�`��]��콆�Y��Y��C�y>�,D�a�z�� ˰$.o�#b	N�r�ɘ�t�ٜj5�x΅ �si���ܪ��Ƴ�d���ܬ�Nzck�k�L5w7��0X�Zu��T�n��b�ηR���"+� i�@#}�͎�I�چ�x��)]G��w���ߑ�]1=�n�P�_
�1~�2ƑN�0Ѫ�g���ȕ��c:#�i��N7�}�������*�4�C�?e��S�Y�V7�?��4�D�����Y����M��p/�ο��L�)�����(u�IIjQw��lh�	4��xw�;���{��'�_���<`�1.��^��H�v���l�;�92W�� �X�aya���i렠���"�i������F���n��g�ix�h91*��M��	t\d[�(�(��=�ɸ���L�R���s�}I>��y� ���R�J��7Џ��A0�����Yv���LpLBi�k���W�D��[�[
7�oT��'���"�����ޜ�Yl8�;�ޛ�w!HRߕ�c��ۛDı��(#ß�93�:��??��Y��;@9�ɉ9�'g"^S�Se�(I�hÿW
�1Dfw���f��<�"ϡ]�]^��H��F���En�!W+����I����~ީ����[Or���oԵ"�(��97���o
{������%�߻�f�]hH�Bd$}� �:>�z݋�=���yC������[r������/������ge���g���zJ��8��5�GO$�zaf!A|�{����uD�OB�C�}νZ�4#�����*F�db!��Zѣi���S�C�7qh<LݡO�0%�g�n_����)u��K��PsZ��RJj���i�<;�@A��KKjn������P4� "k^�����r�Ł�7��߮A4γ]�Ϭ�/&�Pe��n�00�M�T��W�>pY�Vf�������l��ɌW,-	��܉.HRAz��O��LQ|8.��x@�)�+�s�Ӝ�J����Ws�h�D����,��7�.�W=\�e�_v�Dc�:��u��+�S����:��Ce,�/�x�	�_������u�P%�΢�Ĕv�.0�>���{3�r��.�y�5�*�E���f-r�"o�y3=d)�E��E�	�V�Otqa���ãұB'���W�C���K=�(�f7�����R�Fk�v�Lǖ�tj>z*x���a��b{;����-_��ٰKqSI���Rt$K���|�_RTQź%�R����/Kb�'�e������}kv<HM���9
�B��e\��:;�/�Sk$c��J0\��*�p:��?z~�2{$�֚]�[�+�ۈ�Ƨ8�k��%�4�Sb���o-.�C�M��e����\8�Y;G:U������(�hΑoӖ����~W~BJ�@�?�g^/^-�
�}#�Ǡ;H\ĸu�hX�O#��z�Gޑ��^
�O���b+��y��A���"�B�s�)M��7�U���*��!�܋V��������p��������sZ9E!�Q���<R�i6F9��X�>2�'q�������/��'�� ?�g6�t9i�����` "�F��<�Cvv�y)�\����`��Xk�S�/B��v��a3 h�s�OB��ꨅ_:���,��	
Ti��\�qC]U(��S���O���6h��Ԉ=��#)�y9(�g�驘;vA�Ւ�`����r�2��&����p��S�SNN��L�(�y��K�Mxy����ih��.$���8J�Aq�*I��z�����:�2M�-u�-�4]Ω������[�q�PM������_r�r��ƛ�D��!q�y��3�;F�ݲ���Z��u]���p����q���D�0����(Z�;��1>^"[$~w�M��L�u��Vض�Q"�1S�=\N�.FZ��RI&t��:�RR3�LY�x��W��`"����FY���L���H(�mR���ȫȐ����Pw�L���Su\Ln-)��\���.mq=��g����s��=?�z�-��~�v�8Om�el���>�Ĉ��ލ��{�^�G,XRk�.%au��8�*"f�Y�J�3���5Ы� �ŷ�(�[	�\��ㄬ��Y&��6��T�^l���l�l��K�h���^Ю
����F�S0[��O�����`�Ry=��	���Z(��S1\�Ca%������i�_���������3��M��*v>���i��t��jwe"���d+����݅�T���pYq�������ұy3ys��&Fa_{#�ܑ�m���M\x:O��Ǫ��u��D����c��鿚�!nPz}3�؄WUxr��8h�Ͱ)U2��֕���|���Su�,�Dpؤ=r�,Zw��ouy�N�@'�o���}o�yW��A"=�ޛ]8�df0��=0�����{{A������z�ދ=�'�ǁ����!U�T<߾���Xe�����~+n��xd ^��XE�?�8�H!�6�ԝ��MO�a>��F�?~,2���c/zt��)��2�]�WFg*F�zRi�b+^g��i�����,n|���K���jp���9�F��(�6I`�-������g��y:�~�+O�uԳ~]��]BV8H9>=�lz�^uj���7��1p��(����m�P��c$bΰ��'�AEP_�6C�'�{b��d�'é4?N�RΦ�n��N;b1˖��,(�,��tti+lq���G?�6AM�)�G��wH_�-��Õv
��	����ax$�\D��^)q;"�ҧ��a>5�Q��T�l"ҸK�h�,�|tvwi���ŋR$}SH3���Ph;,:��I~���N�-/�`b��0�4�Х0t���h-&��S��A��Յ1S���I��Z�T#۰�����x�1R����=��Ļ�5�,�����!�,��vj�5͘`cl�ݰ�l�*�l����x8F���Y��<bU���5�܈=�:B�Y�����џ���M4~�,	f	��V���
���ϑ����x�D��G�T���G�g'�j���.!T�L�ؤ*�W����b�K���#�����~��=���1�T\qL��gZ/Dh�y{��@Z[�ux��2Y���̀G��Ǻ�,h ��Nw=���복�cӷ8pZ�,	����Q9�zf��wBozp��?�߳`�D���}+{�G`������OB�����y��!0��bL.�fLx�_���~���
�j��J��J�z�C'�d�FJM����;�Lq�P���qp4i��;Z���,k736z���cc�?mx7<
oC��ٕm����p{>�tC207T6��({�O���Ͷ��5m��3����ك��*'�10�>K����zk�E�~ MB���?«����xp�Ռ�8��b��n���&o��)�U�Q	�[�x�i���o�;��G��v]���+\狹G�"��)�_Z-ڞ������b�2��y��4��I�Х��=޸������qJ��f�t��>�I:���Q�֕1G���L���K�B8ߥA1��  t�Sp��������fot�/���������6|���S���aD�Ҕ;����u��g�ӭn��F�w\p�#�|�协�9�y�$���(�����!�t5�Qnf_��}�:��n�����/�ߊo_�p[ˣ�����[v��f�7�6��A�����O1���U=I�޹8t�"	��^Q{2FU��0�|�D�᜵�]>R(��O�����Lp�xn�Z��g���78cFG�<��*�Đ:�1g>E\ӟ��M<^��[�����߾{���
�Oj�z��P3=��X���i�2�>O�&�P�`'��J�G�'�e
�W�p-V#��T�x1÷77���?M��H�"=F3�s�|ʽ��rKz��|*?=f��2UWK�2�_ {?[�F�#���f?q%�]�ތz�<ː���&�%�<�܍��0S�TUĳn�0E/�ݟ��ćκ��k���Q|�L��jԥڲI:�^n&Ý��I^�5"̊.�h�wښ�CY�,�8�?�lz;������B��$%&j�Ag�c�C�����k{!�Q��kET��z��W���9b���N�o���|�+^���G����~�и Jl�SC`R�-���
V�T� �����h�fL��y@���Mp7>l�"	�xQ�|�b*>(��� �)y�.G��dv 3�r]²$��u�XeR��6Iᬣm˕�E�+�M�����j��tP��j��o��J�Ԡjq�a����K�#	<g���	^;&zt⇓�I�}܈&��_+���K����� Ld����M<������k�=��)��nR�Uz�7�����!UC��)���
��_𩖽+(@��yT(��	�J��蚆�Ŭ���ێ�oiF&����⥄lqX������u��������1�2�@�`*��4nYP�w`�?y�_� �9��P����dQ�Y��َ������s��\��͈�:7�4P����wq?Thq'��(�7ͣ�g0m���CCo����+����^�;��!��P��:���#�g�0�'͑����S*�Uѻ? �(�^|�r ��c���MNi(;�u���L~k_)�P��9�9�̵``HD�*��'�a��p�Swy���ߪk��9?~o��D��_�oZ��D�=#m�e�l�I1܅E�Ov!SF���Ao6�|)�kȚ����yIw����u�U,�b=R�����I����˷i�Z,���m؅O��;;7�)'?� �Ӊ'����nwH~�(ˏ����Q�}&%cSNZ��2������ſ!�G� ��?X���m ��d�.��'����Y�I����;G��Xr�N�:~C�a�cN7ŭ�������c�2����i,��&!5�V�9(!E_���mb�G�lK���u_h!�{jYg���N��0�� ���X���k%�r8�Tź2��~�Aʉq�Z��4;㰽�)�]ү,�c*F�yJ ��P:>RK�ME�~�!�Md�*R{b��B���3��'G����|�#4�NTԍ�B/'RQ?Z]�c�=�PY�*�&`��C~>�S2�����oU�-��qvwo���)����G�1�"_0)�5?ԧϦϺD�Xa���7k����K����f.��p�I��5��G������Iэ0�±��/9���F��	� ��v������i�!���J9�a��1�!��)-d))����@���J#��Gl���ê��D���Bw0����@/��x�!��0�#z�lF�i(��xy�·Ҵµiz6=�蔇h(7�?�[1���SH~��0��q��S��� U�x-�i�>��{`{��p���IF��I���`�'f+��Y����q�#�hI X�h�k��M��j��|D{���/�����e�vR{�\���
ʖ�zz�ٖV-��h��E�x���4�%b����x;�}�bD9w�u�؛���401�j�%�,�\"���m8Q��7�&$��"��~��t�O�w�=S"��!�g�)�'U�#D��fo�z%�F�!�M��C�7���ފ�����7c��NdQ������`I�]���,��Pf�`����Jt�,"��QԷ���������J}{s�����g|��\bVIvp��s(F��̖_b��i0�%�S��D�d��B���ف.!�_1TU�+8��� ��F)��pX^B��G�~��&] �\�,Y����%3	`�@�sX����!�;�F��\�h#���_80���!m����͡{��Q�,W�'E��^��wD��r���#�w�Z�S�YtԴf�B d��G���w����o�]�����B��Qq����õ�2OY�7�9-��s�`κS�+8&䷦�bt�)�^�8W.i������N�A�����1�/�+��k)�7dKvs�Sz�>u�=�'������*�p�(�n�8�ށ����-�d��'TX졻]R�\����2B��]A�	C3)X��� �0����E&�Oj�Oyq<�U:1>b���k⌒��ht@�D�� ��'%@��D>(�7u�����(�q1j��9'�Y9��QC���.�>:�TX'�/��Yf{?R�s��}(Zn	�B1��%�o9Zig�DN^�E��~)�`�/ˁ�����&!!C>���y�~��;��d�c�w�-�g:��S5sx-���p�����݇n*�;�:��8�g��@���%�"<��DS�vp��og;��&_�:��F���o���4��g����E�U> ��3��,k��y欪8ܑk=�y:M�5�@K]�l������S��k��؜����Ee#��q�\��$�T���h�T���)ff�Ƅ��Vs���]W��M���ZΜ�'����+v.�\r��'� >�[諸��W��������?,�kb�^n�A�����h4z�w�s�ȉ��ȡ���������Dz*3�R��K6�۸�C���ڄb�0L�9#'>` ����<����m���٤���CƎ��J�E5�7J�;�Ѩ���]?����y��(N�Gz�_�{�`������ߕQn��W����QY��M��Y��e�<��.��g�]���$�i%<�h︯^GwV�s�K������H��c��C�o�u��@���Gﯷ5�$Z�J+U��1Nx:��Z3Ĕ� GE�7�JKe��}�i o�,�X�I���;=aH�Ѿ��e�(,Ǡc:��%����^�>>z���:����<�����7���D�P�y�N����%Α�SJ#���\wV9����1V3c���EE�N83P�Z@+�[�Nc�	�����6ínIY��niu'-k�`���q��	(����&��9�Sx�X={��o������C���1�̙�u�?�3=;�����f���x�ͭ�df	;߫շ��A�|�iVw�7��M��5܄���r���������h1iy�N�Ȓ��WU�R�(�nt��^��q�ѵm�t��B��
��6ߋ-�����$��ٷ���g@��r0�|V!�T�V=M��Rj�Ҏ�'v+� ����_2zX_)9�٢�k��y�3T3E��:I2���;�W������1��WL��I��M��E�C':(W������dg�<����u���fv�
ZX�۴�R�V��ǹ����"�sL�v��kN���y\^�a�9M$-��?N���C���� �r nY���dl�M��"L~�<������k�R����r��=�SVz��>A���ݽ��FP��p�)�+XgP��{�g�ā;&0 � ����\fi�R�{
ѐjke<Ӡ���� �<
�2���t*�QNcx~e 򋏱���T>����N�|���x��A�߰��q��>w!퓭�ug�*���)��;ʲ���oӸ#��;塔��@H��h#��]�|6K"O`�yߏ?�4�oL�&�U�6�p���$�J��-�H�����P�Օ��<[�F�in(�H~v��K���-�%���,4������!H��.���K;�gE%z'�l悆dyN[�=Yl��Φޢ�4ٺ�[c������n��e:"g�DQ���?V���7/2k�*��Y;�2bTA����c������R0$�4��'�R��"'|�&�{����Z���O7F��㾥�lE���F����6�cW���SPs�E�3�Ze�/>FoޜP�d�U�l��<w �c?�T>h���ud&�Ï��T��r�	Y+\��_��ͥ3?_�qf��GE�kX�A�Z[��'�?W.q�F���e_e���<�1sӚ�΁ؑ\Q�r.�԰%�s�I�i���9��탼�e�$�!�г�Z��R����X(�s�j�E��z����5iv��ȇ4j5��͗9��Q���/�-gf�^X�}ϛ���>�
�T�m�}L\���?M�'�$��#j���lw�tqҸ:�Z�_"��Zצ�Lfƴ���ܨ�L�����~�~`������[^�U�cL�߫R軻��#�B�;#�Xh�d8^͍}Ց������5�Na����$�Vh�	�9����ꖢDJ�f�#H^�qXn�ts�E����=NPɽIh�Ƹ��}��Q
�?���#����V��{�K,*
y��ӂz7��;<�{-*���$��a��=/�MOǹd�/U���?����Xq]�6r�ֺtH��������NI��y��K��E�j��р�/�n
E�jcY��瓔C�]|�h��?����&d ��&�/
�������}��֖M�=oʎ)��-��	>���z|�����pMe�b�pI�,3�7�:���v�6�r�`)-�Bƀ��qv��x*l���&3`�����?/	�(�{2w���'Oӳ��Ƈy��SJ̑PW��7ͱ�M�OJ(���j\N赝��>^9���G�ɼ���]֮���f�K��w���唕1������}䜡#/����������k��#ˣ%غf?1{n��حDu
��D�.-V�%�.(�%-v�ċs�j�j;�;ǚ�If1��B��G����(����(r�v-Ktd������f!��6�P��w�+�5T;O�RW��������
�����a2nj�2���q7��Ie�㎧�YV���j�YO�2���� �xt@2�Gӛ�_~ܿ������,�#9o�zBx㧗��Q��R��C6�n���ټ%�>_��ܽv�N��_�7�f��ױ ��!LQ3�B4��{	��3zޝX~;Ѭ�m���f�t=T��)5d;�c"~+�қ�S+(��C�f*\یj|��E}�Aw#2�Ka���D	HJTc��o�%P��Q���\��?Jm��dݠ��(g�{4G�%��M�pM�
;���m�w����RX�2�.�(1q��d}8�d��5�a�Z����{��-��<���Ɂ�������w �`k��5
����OCe�]����"�εJEY���k�z9HV��pF�CK[ >�gy=�Ԇ~ܪ�	}�*��s�C�OK��{�J��}�����uwaw��v*0�2��=��3���z��S<��(���i/Ƈx�����rr䓩P{���J�Ӓ����5[��+w�5>��`�j�n Z?�Z$L%�8���z���GbIw�rc(/��R܇�Sz���=���-����7�� �@��N����Pn����zVCo/ar�/8����Ƃ��T�����H���t�̒	u��lN`2Igm!������ZAJ8kb���8�߶�����u�afLF@��߯�<���n(�Y�w����<���D�	�ܐ�׎�?Y��w%�""��弐�O�+d����sf�nI!���NrV2���9��9\�Ta\��5n�*�X���q��-4�8<���p�6���q*���)%c�kj��k�����L�a-�������-�VP%zs�_�CA"ó0�&���D� �I�u^�a�/5��c�b�u��xj�bR��[P��űۄD�mJ	9�5�L��L��/�͛/��NT��g�cNn���s�u�cx��oVov��
�2�6�>�$�a���tX�b��o�ٖN6�?a��7�F���?�8�6_"B<�b��9�x��RA[U�0;7��fwW�E��Y��z�Twŵ��S�]L!g�̀�0W�l�c!���ōZ%�P:pɾ������un�~]W���ECS/�B�����M/��y�	>di�w����~�]�af^��Tz7B�}��ϸ6^��g~�J�J�����D�^%�����^�{7�U�j0�Bp��Df���J ~���`�"�L��g�SJ
��R����(���5�``��lF>3��򩒳2�u���X��C��EX,����N
��b2���y�4��\6q���%7hps�\��K3*��2��ۓ*�H��R��V�p��r]�Ωo��/Z�~�Ҡ*e
f�p��ME¼P��Ԫw���>=�s�˃�G	���B�j%�vȮ�IĿ��҃��r��=\I]� �`z�-�XI�g���������DCbE$`2�&#��������poi:���F�i]xX��[5���W,�X���͇�҃S��|�S|v��.X��g�d��	s��E�]�Գ������M��C:�?�~:�%j���ɦ��7�L31�u�g�%������V��!��US�E��Z�Y.2�׻]��2Z��5s�G���Z��z�H��8�����{�ײ��Ϫ2�ʌS�T#xɼ(
�3X�.�s�^�0#�~3�>r&"u�8k��(�Q48�랧���8�l��'vr_��?��j��^�>]�W�����1��%���� �s|��!q�L�il���)]�7X9�Av4�١�ܻVb�i�0#5��Y�X>y K�:�C�L`ll��%�5g�]"6H�L$q�Mتظ��d�*y?ڠG;�048���v�Kb�$o��f_�@*W��.�����rjY��7Fţ����a���]�U��H�K|�z�����;������f �P�����b�;)�ە��βC����FwZ��`K�?uj@��\���\��Qzl��Lp��4��*�GK!������7D��7	e���pD��4�G?��c\��ɍL�H����6��}㲜��_-U�gw���؁���A��/Z�O#�����g��~"��[�ڄj)���5+��vk����Q#f�ؔ��{$�H���Z�U՞���>�_��>�\�u~��s^�q���?���b/�aP��)2`��]���	]hZ��}r6���!i����W�$�	�}\z��8\��Vtj�"�I����j�<�����x��4�9�.�Q���&��o��Cw��^�Ҝ8�
�.Q]h�H#q�N�<4.?�:���R�����h�b�\J�ᗑ��m�帐��:梨�_��}i�_-c�yk%�i{��c��=�̏_X�����gGg��u�E�-��aV�=9�"����<����&��W�^�m���\Y(ة]�Y�D2)]$c��i<���(�0h�6�3N��4��]�z(���8�Ӏ>��ً�vw���F)�'�<�Q��/��5y��=W�?��
'�Lo��y�#�#�%�4�c>����NR-��_}�e��m�kJ�����	K��AX����2o'�+e�%���|/��Y>�dnP�����]#7��l��/Q�a��#GԜ�������P�j�{�M��2����%St<�(��v~�nԤzx~]}̕�nNk�h�x�|��Ĕ$����.X<�i|��CE<@�X2(�8y�Q�)
�A�CӁ+A�BP�S8J0Q]�j��W.ՃP�߲�������ӛ̿)�t�y�Yl!_�EW�?fiw��Lu��<Orr�'���x��ዯ|���{��H�����n�H�ȩN*�����D�'H�^q7jI ���G�I�c�r�y-���Y�)am�VFj�=Y=��)+�_޹'D�������&�����о[?�|Ru]��G��~?*#��Y�z[�|:Ef�ۨE����F�ڐY�JNQE��}�RbK�OV2
�K��`֧�Y(��!`9���<��|=�^�=r��=&f�2P¡�tw��
�!���S��=�
w8qd����d�C���4�	R�Tr�����G���Px�&[�R��C���k�n�yc{N	 ��0Pi���ys�U�f����5g�e�i� �Wej��M�b�nm[�.��]Fp�e�W|�O?�?2�#A5�7�T_'� �c%�>j����O<(	R�Y��G�������@2b\���7:c8<�ֶ���^wd=z�h�=�0�y|�}��M ���Z�3��o���ߜ/{csNx�TĊ�]p��ʇS�UF*��S�͉�Q�H���� S��lM~
���L��q��n̿�b�$!'���B�I���ua$���NՓ��$>~� !���,Qt�׵4Ț��,0�6:�����7�l�l�a8d4��IW�Wa�ޫ����gl�x.qwi���f"�/9��ځ=$�k��E��.�`�۪��RP����u$?L+-�h������aC�ó�j?���)��k��S��D	/Z`�����*��[��xv�ˇ�f�gt^��/<�������jֳ p�E���١f�ܮΔn�����~]	'f7W��i��jl?9ݔ�eOm^sb�s�F�r���)��f�D[���v����u]F�o�kx��I�%������vf`�rS������(8n5�W��R�\I��4�@*�w�k�`Q���ZZ��mV��d��bXb����AVgź��	����nCw꽆ƒ�=_{�L��w-5��oc����$��|l���t��e�5�l{Yb�F��V#m@-	�����e��� ��W1�mG/�':cwgg,;�j�j^�vw����ѣ�{<%�����B�
Ύ�k/Z<��pjʖ�m߿E�>��OI \��3,;�3q ��Z�#���<�q��N�LU|�rh�� g��3Pgg��F4����$����0����`eP�8�l2�1TY�T�'>"�Ӎ$l�}lY�"����~`��� ,�P����m��:M)���#����nT�b���K�7���o��F����E�H۠���Z���rJ#�j�n7Q:nc+:��o�[�_����}Q����*n�{HU
�����U"FE�Z	+��n�+A��Cq�Py8�4��xeXJ1�?�X�&S��XQ� -��ʩ�;�� �Vm��Z��� "��a)Q(�巴���N���㯒@���o
]"?��R�Iù�'?��1����*�H/Q#@[��a�P�̮�|����f7�A?J�$�#Q�{��K���m�b����~��D�9��<�o���5pb�O9�87��r�^!���|��ٿT<�+]�_YCVj��2߄�4�Sݠ���M�ଞt�Tp%p�'�?��L^O��萪y9u%�AW�
׳��!Р����3`MK��I��*k����)�-�(L��S5by.�����|:��2;�1���l�\�^���/w>E�6~��׼egg�e�>T4Liv��ľ�wo����o���W2<�I�)�G�66j�(�q�^ڦ�<+yU�^�̤5	���௎L�)�W a�p)���䧯)������ry�>E�!ز������W�a}�8Y&���@��X�jR�u��Vm�g[����^+��)���:�S�i�+n-|�A6���u�?#�4�VvD|���(�6�R�HF��3$x���3$�r�43y�>��m��y�V����I�I^W��*�ٌ�#��>i�d����������غ�Z��NaS:�EIV�6�-�
'4���E~lp{:<-^�?#���~LTet�n����B�5��ab�@<t9��F`xdr�w�"yU&��S�M�=�<���yP��p��f^���B��\�7�^r���t ��G|�����=��t��LBA1�R#v 5������cu^}�kZ��|,ׁ�&�р�!Y���ׁ,�w<cXP,�r�y:��%2��,��7��_�XM`����Sn�c�G�]�ANa%�LG���i��}ΛzJMż��g���)FXOTg�͋�#���aX)�����������pW*�J@��ʭ�,�H���}��B��a�|ɩ��R!O�Mpw�t�
�,�e�b\U�A�BW���XM"������:i"�;�TGE&fM�oǿ��Q{Z�e�}�GD�@x��K�6?l;֏����܉i�i�6ҁG�]��w��%����w-�4�T���[ tb�:.5�q�ba�1�Oi�T�;W��4�iG���U6e�=z�4_
v&1-k���Z����j?G���Ta�2��.?��}^�d#�?�G�Uʅ��:�]g-��اS�W(\\4j�c�AK����`� �9<�]-byv��VH�2l��$�Y��]�<	f�@�ɜ��o�_;-:U��VY�<� _�1�-<�T#���F����c�&	@�^���%�����훝$o5b�����u�r�:�{�"\('���/��3�z&��{�����/&itci2K�·j^>�7٣��rF��^���R�Ø��ʕ���+}�����L�'���;
�A�"  �Sk!�Ӎ\ l,��d}᫪n#���p�a����y��K��0Aʜ(��6Z�Wl'G?���9�e����箟�w�M;��Q� 0�y��.Z(-Ow�x5��m�Z<�2�Y��[� "�4I�:hh�y>m��"z�)���	��8c���� 6$������{���SN�ώ[�W�1#M�������d��{�z��_�l�H����:Q�/5�/�]cټ�|��В���� J���.;͢�'s�����D.AsNf*g�Z^Y��>C�����Y��{�u|b W�S���S�x�,���۔pnÍȊ��uTD	/���b�3��oX9�>P��5%1w���>@]{��`�q����τ���ڏ4oi���̂n��a�^V��߇]���6�u��sI���%�a�ڀ��X#2���iO���� �=h��[q�Cy��n r�m
sceQ��4��j�M[�	��m�*x���:�њ�p
Y�G����Q<��Ym��׾&MɎ�	��5��E���#�?s*�]�>���eqn��+o�{f��b�ג�D`��a taqt��XI%�X�w	���>�	����{�P�� /�p��&�ۨA���'�xQ���f}m4*>�����\�� �~N�Cc��N���@���D�h����/����C��D&�x 𽇣f�;����vaշy��N��
��3����?�����Z���h�߱��E:�	� �+�^I�y�Z��<u�:*�zN�o����`��P�&��������� ?4(�?��&.�-[����E0A����!���hګ���#rےT�!��}�x��I�-i���,�9����%�8�P.�28����TM8�c��Lc�Z�<���%��Fm,\9��L3CYѾ�ۺh��%��u
 ��aSD�R0��=�֍q�m;�u"5�K�)<��]G���c��s��^~�yL���KS���K�9�&-Wct�&�[J:��Q/�����s3V��}����/�pufJ��h�7+����%�-������8FM���mG��K)�@s��6��_vZ@�u����T�d"�҉WE���y>��4ˣ$�'�I������'���h}�ج K��Χ/r~u��gmz@�hZb1Fc�y*N�@�z������`I��f��Ͳ�������xbt=�nB	v�?�h;�8�:ꢋ,f��W���x1ͧ�эJW�[�c��}��r~��3hRd�}�5�����ՑCE����x�K4ز�n���-�����*�H��Jm;ү!�L�3 �[�O3"m_{*��-�nc���?e���������(?�Z�e$�#�lpu�
�����8�ψΙ~�	
]��ԕ�φ����d7�ox�X���e��6�s�1�G�1��RMN�`^_�V:op �is��������+E���NT��	RC˿��|����V))>�����)S�����^�j�3���]B\����IdP������o14�|�tS1��QN�j��IC��Lb-���۫�][\��h�����Qki��J����,2��[�#��a'��z"�Q�Eܔ�
�c�tx5�sW�j
�yU����U6��X�B��$`F^ś��&QE�@�;-Ԁ�\T:P��� �~�n�-tGd���d�H�QH_��t��r�7V=R�U��w+��5�4^�.r�����}b��:�&7��p���v7%g��1&���5���U��^q�E<M��e�{�K*�����\�7��*�(��c�.��ex32kv��`�{I��� P�fh��,1_�z�2:�d4�W~���3�m�o��ї��ܗ ���\��;�vc Ӿ�}䬋��)矜��/=$ޥ���d
��A��z�n���L*��QqD�ݘ���(�����toi(3��.z��`�݃rqo���3G�?H��W!Ƭ/��T��T�zkoI���%�)A��zN/1���l��BT�n�H�A���9�T�rF�<>d�o[T�g�@��gR���,�sJ	{=ߠ��]:6/e��z�L���xt�ٰ̗��W���E�DcPeO_ȕ����O�'mHMH$�+u�\�����F�!�֯�2[��������YT�J-'�x�Zu�*��U1��s�g�-��3M
�L+�)��eӕ���}��:��s���D�S��������*�I�z2KM��edR�\H�@s��UP�G����yӳ��SH�M9��pH����b�TV�m����!�`����n��*y��^]4�>��e���R��ý���$e�ޝ�#�弦����� h%�,�5i�ͺ���|��Uh�� �g���*�Ð�Bɡ7�'����#�� S�0�n��Ϣ�ؓ���d5�2߅��I7��F-  �w�/�� �c�7�t�� �,�5`�O7�w���EYw�~�%��H�b[���$�g�@Z�y T�>���@�n�,��B�&Ij���j���`�?Q�Q���9G��.:�O?�i)�z��>���&���	+���<m�����r'&��N�S��q,9���`U����ݷ�}="����w����Y�]��m'�q�A@���\�I~ݯ?V��ܨ�{WM0�)S��|C�q����<���� hu��b���J׭+�ϟ��2���n�)�K2��/o�5i���.X�'�ǮF��җ��#��3Efy�rG/�t汛K�ŭ�鞬1������ey���}���D�f#���V�S�w#
Y1Zn�����H�vN��K	�`����1��}?�an��2g�q�Y,�:�fR�$5���bI�'|�o�ةU(�`�]��̽�����;�z�;��h}9�^vc�U�L���E��< rq~�=1f'�?��h�Ke��L�	2	�y�@����
;����Xg����,�`�紣ţ�'�?���9���Sk�6�@`Nӡ��i�Z�b� ��Ӎ2��~�ka�닺W&�=#��p��>��X4ڠCs������}�q�g���A�-�A]J�s�	י��I��mT@�vG��AX�/���8����`�\e�/�PG
y�+4)T���8�}�_F��y=��Ы������4y1��=൷���T�R���__j=ų\��@�Y G�<ި�,��`R5��[���������u�S��d�S{�p� �mŴ�N�����l\l�7��1A3sq�cD��g��ajj&k{"�S܀K� 2e1&	p���g`՘����R������W��쳛:����8��π�՟Z� �< �9����mJ�ϧ�\a�K��A�p��0c�`���E[�~3߇���������
GX'��|�*�D����150�R��1���Jp�G�H���7P�~��֫Q_;a�|I�T�L��X���Q��ަ�-�H����rsŃL�{�n׋�%�"�{�'*T"��6F{WCorI��LϩRl�M(� �3ݲ���;AЂ��/�����L��T�;�`�o�7� �m��Uz��lD�q��Q�Id�AE�`��#�S�W<?2�%��|��~�N�nh�zD�sc�@�r���?�1`�8U��w: i:lEU���+k�����>�i�4�;����bMT/!�D�޷�������^<2]��[�FY�^2{���~��
�ئ:2��*,�)��oly{���$y��^�:`�`n����	���.�����F�_?�[!�M��0����ލ�2�(T~�w�iԺ��m��E,d·Ap?aO�:��~�|��>,��΀�	#L�����.*��No�p�����s#tR�R)���q��q�����[#�अJ��s�����.�$���g�<%�Vk|M7߿�˪�N_�|$�K���߱M�-2�W�B$AМ�3l����+�t���8��������"3`
�+)f`���!T�6t�66�"����=y�[�ܶ�\�M��hR4� ���9�J�Ip�h���9�6��޽��'U\�47�B����#*
5�C��#H���1���#)]��'{����Q�Ф��k�[�O#��-�pp�,����k%$v�:��K�~�w�Zn���k��~�E�m.=�̓�=O/���Cxa͂��z�}�Bo6�&4�#W H�q�ߵ}�?�W� ����6ڟ/jmg�]q����fd=c{��:]ͯ��|p�F� �D\�B�N9Koxp3�t�(v�-c���ȇNA�Q�m�N-e������o� ������ח�3���K���� X���q���1��0)�n��߾ᡕ3���2����"P�m{����+6`������� 	���ڬ��zQ
�h(�0��"��>(��βn��|#~���z���7��^����-�j��1�������۽��>����"�;ܕA��`K\]�!U������M��b8��"�	�d0�*XB2.��ژ�&�)��#<T�_���8�߻Qm�ەt#LP���;0A�Q���A����L�=\�M�!V���i8ѣ�8	�4�E�Tf@��Z�p�7����c��i+ah$QgϜ� ��:4c�8r(���vA�~&`��j��(@Ԉ���m��f<��F ��j�kY�6�|�e��B���}���I�oP6��X��z���-��m���a"q�h���[��u&j�{����4_v��J�?�)�8���xA��W���e_�.�Z�iK�C��^)�M�����5*���-���.���w}! � x~�������݈��<D.�;��i	+2�h�Ͼ*���#�^c3մ�&����w����Gb��%Qk穩�%!z��-4X�θ�/ �9jqt��\��4x��y�}��c�VĝZ��O����^��@��u�_���Z?��H�-X����w��E�6�ߔ�l6�����(� �9Y�j"�>��Q�z���(F!�O�u/����ط��=r��V��W��BP�	C�(פ&�XmBNi4��"r�I�w����.��~�9�%=V*׼��n��\Ey�^��eN�3��̳en�߹"aE�5���g�C�l�_\��P�a��+�=v
P����f�?���d�f�ë�=a��Di���2b�j�2hSϢ��:r\(ZGä�P���ȒY@שAcDsxh����.*�C��c�)C�U;8�f_C��UO��+�#�3��BS�%��c�^������dU��\N�/�X��}��K��ٽ�RM��ֿ_:#;1m�6�(r��y�'�����'x�q���ac5V��r.�U��재"4D:Q�%�l�;���[F���+m�v�d	wI��Ȅ��k���J0��_vlK$K�e0�Fi��63���O�\_B�`���k��Z�	߀y���K[N����=�:��k'�vuQD�|��u�_0[�m�'t�yw���G��|^��$H�9>� �$�
!�w��<�K`{�.0���h�o��:�E ��JH�1���	N�^3�s�M�=<��Jٌ�m�����x�&� zRL�i��h��y���c�������F<1�`D`��F���_R���^�-�~=vC_SzW�$eG�*;%���=��[���X6�۲�\�ID����?7YE	�u8��@]��_Ob^#1r�����ݿ��1�
v����U�V��E�>��>�ĂZ�d�O�����~e����T ��3e��W�2���h��qq�g���ݝB�32Y� ��.�w�/���+&&7�!�)�_�;�M<+�T702����
Oc��OӾ�넖����ބZ�~��,&P!G��ۨʁ�����9�&9~� VbLT��f@���p�YuN��5p��l�Ek����i�@`��.O��]2�UX1��Nbv]=� �U�~��Zb����̜��m4m�c�/IDK_� P=�F���#'��;ۯ���7�-����S���,�Շ縗ńS�4�wԚ����G�ҶGj�$��Yk���b��P��(��N�|\�<��3�;ZO�U;iW��2.3aFF�����(KC��e>�ݜ2�^��(w!����:�D׶UF4���h�tx�hy�%��n�/,�ɔ5D~�{�)w���~�������4|������$��tUm�^Ջ�z�맷�>B��"-����<8��9�)PL�\@��rnDk1::�pjȀ�{^��A�URD�߇?��p�>y� Տ�ܶ8�����
��%��Y���kR�������S�*.�3K	�MqD�s{�A�)-g� xg��_Ap+�N
�zQm�y�t�7����Hsb>����6��O�<�f�}0���
���� }LXb� ������[�Z��S��u�g�֋�Rg� (���dI��3�-���-�0��N�� X��s�i@�,@<w�p��\���ԃ���y K�Se4�V�]��׬n���84���B, T,�1�E�^d���u���L������D���.b4͠�V� ���r�-m�;g^��>�핱Ϣ�L�v\��]t�I-k�|��T� S�����m�t]���^�� R��\F���̀���6�~�H��St# Jzʯ�'�4^/����zw�6`w�߶1lT�	%S�78�-J������_-S;+($�_5r�;{ƿ�=�d�JZ�2�O���7����_p\��BS�E�u�&fUlv���ya�=��9t0����xXR�䑒?�MȍjҺl�_�k�#+�jNr������:rH���J(/C���������3w�n\�1��#@�7��BG}P�<4�3�S��\��=@F�49SoBv����>��X��В[-���mX}���i@��d�9m�6������* ��
��ĵ�>ĭ�6����3�1����Kf�L�Hp(�^Qv@�G7�q
�Z��C����_���K�M���[ey�v%�h}]���Ks�i�z��s�\kqa��M��E:�� n%�Sd�J�۶�.ށ������=g%�W��o�b[�#_�ޒk����U�n_�~��#��5x�J
�_D>EP�ڶ��E����Iv�q�\�ك�c�K ���-|� c� ��9a@Ob����=ñ�Lmɳi�_�z|��p�lJ��z|��׎!��Z7r�n�Y�R/��>^BQ�o��)��\d��!�r�Şm͓�j~lu\]��̀���*]�����?����+��iN׋?��E@1BN�K����V���|�$k�4�x���?R���~��-͝��otd�����=,�!<��6�[*t� ���]J�8�����,SE)�Z��4���v"��0V͛�*�(�?����o���5~�M�=u��x���ɀ��vI-���8J��LQ���J�7C<(�ʁ2�J�I�,����'^܁�X�yI��Y�q  �h?S�[��f��rM�"�%�mXb[ݓ�av���ȽS�@Pn'\jd����n�5:�ؼ��U+��$^i�~�"��~�dn�8u&}��!��w��`kk��d$4#�ǀ@Fk�09� ���У��	�s��C����Қ�W>o^���E c�$U�8��v7v������~�}���k���a�]�Jݯo��S<���i�5��Sk����?�A�,p���g�eR�S����I�6yuA�hxr^OLw7`j��'�F���MA
�s��c,���Q�i�S�3�K����6��:��2��H��_�����+���j��Hu���������A"ڡ�E�V��L1������<5�/����K��cE�mhh�v� �$�Z�nFc���Z������8�E���ޚ��)~F\�X�<�m_%*]4���2����'�$�:��\a,X%�؟��I�(+��E��S"EJl�y����*	{2':@D؍�o��Zѩ�ڛ<����O
t�J�8��L�{0�z�qƜ��E[���}��I{��@�ɷ����76�;��TWZ�_���zR�{)#f�(�x�+����K�<@[=���\PW�YOm���*\^ �~$ �yj��ȐRb�y�����8�ݣpS�E���6��Ug��4�6a�đ6��7�ƼT���ڒ�V}2�o�9�����l���|�zp�'��B�e����
��݅Er&h#U}T��I��:��u���9�3�B����7(�5&�(��ǆѰ���Fr�m>�4��,=i��}9-u��_[�	hXʥW)��.���������Y3k* � ��������4k�_�u�-}�}L� P�i�D�޻��U'�_�I1\��%]0��履
�>�����w2�@�L�eQ@!xD�֣���X�_��������vrq�{�����JQ9��P����/��6J��f�@=j��� I�.4�	�tL��a���(/�x�w�(�9,4��F�,�z���Iq����k{��1
�@�j{�>"�h��*5j��@���!�-c�A�7���<��}v����&�v����Ro�r��K*�}�E�4i0��~�Xk�A�M袝�gE������v�w�ޮ
9�<�r�/E�RH�f:.����-�NF�[	��-x��Jͱ^��­�	���2����æ�1�b8��f��x�8�ǮU��ʯƘ�>n�6�UW�Υ\�)����r���]��^?���jR�;A�� [�ׇ��@�"ľ�=�!���n�HXWb��~��\�����.� 9]\]�����y��A-�1=���]�3������c~C���$����1*���@)Qͫ�ϕ��ͳ�O����߽�8�����Y�!9jy��S;~�$����q6��j#�ͦ�	只�à�"�'7���e�퍏�XE�@C�1�:�{�p?�HUv�پ-V�A-�3�K l��t�g#������(��	��| �/�0Ւj��8���~:_���ǄP~�g��y#��kj:�Դ�ȃǻ�4�R���L�eڧ\j�;%�8����lǥ�
 p��G��؋7ɞ�b�旸L� �-i0��k�s�p�ݷ��D�m=Nӆ�Oܢ��������T����'���[ ����Y�1������ '�=H*�Vs�U��B耺[�s]¹�TT@��Y(�ӭBEtƏ�Tp�lj-&��F�Z72P���z�D�&�f>�������c ����O	�/2�-���W��>d��! j~�sb��V���R�<��?$�	�ٔt��Fr����M�� $TZ�S�a�+�Vp�E�{�|cޒ������O�*�,+"��(ߠf~2M 8�Fv�<��g�t��.�_2�	�J�I�N���Œ�`񨘘����8��F���'��1�;�e(����6�u�'!�tWV��q�7-o\�X#�w����S"��?pԉ4"Q!a*��-n��AS�Kb�02�v����뗆a�'���{���}'���-�ؔ2�~�kg��cO�ye���C�7��+ab�I���X����6��$���1r���E=�~���$"41�J'�D�Q?_��'�l p��T�y��u�����7b���n��]ѱMa�3͇S�36� 5L{$�$2S烓{l<΂�ow��x�5�+B	,8�y�_Yp�_'sro�vw��ɖI�=}K�;��|(X�� M���ӑ��pIx*�����k�g����ǾIgd\_�=�m�8�e��>Β4�;-�?1���"��DR�_�,L�}H�S@�~�<P��D1��@M�J�o�P	2�P�e���~������]��#�2�H�G���r���&���S�|�p�!�j�zr�T!c�wў�3�N3����/�����\�E���q̫FA��+�?u>����s�?��]�Noϱa+��*�6��͡�",W��+����0�Л^�Ե�>��_�F#���]�e�(__ܭ�z��:'�WQ�?��fC�G�j�)�E�Y�V�n�b�~�p�Ca�_�=�hm1Fewz���׉P�c�K��;���dV�G|�[���r�/�[�� 7��\�e�Ԓ��֓���y�`DO��3��bp̌bIfG5c�	Y�k�(E}����;�K����!f��l��/.� L�o3Q������$��;�ܮ��NZzhwJ�]q[�Y�lX]��ClG��`��јƕ9�sT� J�� �����k��ʆ~Q�BOp-�FHP���%�#��"��j~w©���W����'���l�&u�qCR��î������ �AY�����bIW��QM��[�G|�#�{;\�+2V�e�a��.�x�ā��@���e��m�����|�-㍌�:�/���YK�P�,bW����>1Dw���}4z0#������C(�YG,����Y������B�pֻn]4�����r!~䳰���c2̧�
	�6*�a�J�e����7P%ܶ+�Kc1����5���%����%�k��Tbi�	� �+bj�?}=q8���۽|�q��w��4U���۾Y*5�fQ���9����Iӂz4���2hG�:xF'/$����Z���U����$b'g*g���>��d��$D��@j�ќ4g�i-}��4��_���H#���A�zN�Y�&"��S�j�K��eX8j��:��|^H���͢��Kɕ��d{ `�s���!�+��o�i�¹�OC�k*��Pݮ�Re���CT���s�S�3�)��ɾ�4xu��eZ��� ⿋��!�͛��䠄�m��(A��.j�gD�ern�2 A�6�<l�R��.P�����2��Ɔ]R��<=��K,:��
�;����Q�=y ��6k�DI�x?DbPx��,�%D9\�&4;�b?�@e�R�����m�|At" ^�԰*��v>�1���K%$=�n��~넨�m+�tG�*O��T�u ��k�z<��y=����*s�K�;���z�%��2>?�i2r؄h����`rx�-�'/ƚmt�E�f�5i^���Ȯ#��PYwu?4��~s�zP��Nċ��dh(Y�37�-�Xo��!�����^��V,5Q�,��y缯ɑ��D�С���g������ء�A�Y�,��b`�~��{Xm_)�����hgDX��SX�dُN�..?�b��d0Y�p����(�#hu�XO9= A�r�P�!�`_�ԩ��e��z��u��u�!i�'��12Դ6(9fA����3T�w�����,0�\�y4��9���2���0Yϓ�������Y�]���Q)������|ͱ�k���Z�U.�5���x�&s�FV>�5i}�Ս�J2�ʛ�s�~�b̿�(�We�G�6 I�ٙ� )���T1"7�����v���F���y��o�F���<�òP�.~�y-2f�y�  �z t=�Hǹ�YE;���"t��$�|_,;�Z�11L�Fp��[��-'�c]��&JpRω�cL��k��"d	���o��x��~N܈�_�c#�����EN�*���4��������%h�2��Ex��5��$�+��J��ʧ�~���ʧ��N�s�� &��{I|D%Ի���������d��,)V��u��D��r�X�E|
 ��y��ɿy�`5P 5����JN{c�����p������H�p�{Y��ba�Ѭ�Cm�t(R�~<s
p ��ց3�a�^��J�9�S�B���ĦV}�lJ�˦Py�*O��~�s�H��*�V]1Ib7pc~6�������7���uP�|�P�<�k��>�V	,�>!C mol�!4ȔE��n��`��1D��30��{��6ߤ~^�7�H����S�&mn|�0"��mau�M��.;�j�T��s�ug�8�&\%"���B|:��hhw��s+iK�ЗfL�*]�9gA��2�zR�i�lm�"Ϯ �#
r���'/FJ\tB<hn9���3T�J� ��.�A
�G2A$��ՐӅ����ʛ��%' ��+Eb�b<"5.�C�������k�}U�O�c� 	�ܭ��ښv\��?.�_�p ������M����*���������u��W,lB�gqs��R"*E���MIU����E5u�o)�A\`�/?���V�NGJo�����Wq��9 �x�,�/���ِ�e�&F�̠��5�7�Υ����O�d04���[(�S����G��l��K���� �aw^+p'���d%��T ��M4\��p8f��3�����=q��1Ę�9�_���߬H�
��ʵ�N�3¨����t-����$���|,��3���0�UӚ?4ǔyQ	p��j���k����I\r�ˏ���]���[œ�����mJ/|��TPg����O���GN����+�ƚF��㼗�@��,A<�y���2H�,�,M�,5�q��r9�\F�wFXӐj׳{#��Os�ј���	b�0$���)��Yz}%������t������O�b!�Mж��{���>X��/ֳ�wl��W�/�]}}4Õ�w4�;;c��s���?l�_\��z�M�8x��3�?@�l�8�`�:�oQ
`0�^��:$t��q�:d���MJ�(�5���tY���o~ ��qT�ذH�#&&��i	��^�;�#.;�d��	�{n�k��_�ɣ����/R��K�����4��ˮ������-�屯�'�\|�q�V\4&�p�Kt���5ԛ�l�ų�[�#Ξ���5>�4E�~✚��2:5}�m������o��9��q��������잷wYXji�i��ZBr)i���EP@I�%XB���XP)i$W:����������3��5����I^B�WJ�	/�_m+�L�u|3ry����+5/V����_>jC�W
����_�7�.�Xe=Wv�����T9x�å�$.��ڟȧ���y"gtKO���%4����dl���@�t>Q���S^WZ#Ƨ���ă��F�R�}���z���k��>�-@s��/�vU��[��3�����p��L�},���	����~�r�@R�\������_(�KU�4����u&2I�a��k����{c����+0�G�/<g���*WQc�n��t<�CKX���U�=z����W�Ȭ�M���O�F	b��w��ʓoת
T��G���W�}ߧ0�&僧�e�����jH�z�\����9���.C�/�rY���#ޘ�:�_�'o�9��W�_$��%�˲�� !���f�Z��P������d��s��W�����7	H\��Y�>����\㏃��_��ħ<\W2é��=��b|bʐ�lH|�Ҷ�M��k0>�n�����◩��ӈ��rZ����s�ӝ�b�`��a_�m����z�!,	���K��x�cѝ��� ���.OL�:C�bG�����Sq6���j,1s��k�^)�*P\���Ϸ�c�:�@��'����o���_�� �~��lԧ^K�vM�U�ȑ�;M<Si�6(�X���^e���*h)<G�痾�=u5��s� #��x����O2�R�?�AtZTZ16D'+
�V��l����C�R�L��Z��������7&��I�><�$^K��i.0-�9��[�L�̋�Q���\/ۤ�Φ'Kl��`&΋��r{=�#��9o!�\֚،<�☣eD�ZZ�H��y�.�\�U�ɷhhg:��[�e~��r��\@��>��	R��ϳ����u(E>�1��^�V���T��DyPUc�B��%��ţ�*4�Fx�'�
���Q��Q��h{R	Q�w	̐�����%���ؙ��D<���l���x��EA�{��X�P��}|�����Ԡ�,�m� Z�K���v�ͳ�fK��ߞ(�B��0�K��6N��r���A\���m�_Ɯ	��H�=�R�K<�%"!��[��_��r/k��׸��-X�ω;�'@8�����H���XȽ.�ǈ����4p�J%��Z���ʤ�c��o��xC���\�>���Z��*J��8���(�.g�l�Θ��pa�u��n�1��EeA����[m��RB'���q���w]��k��u�
�
;���#����#��~D��Q�
(��U�>B��dbN��=�h�؉���eP �W;�5�w9��ɺx02�}�b7�^���O| �|m��$����dnr
��ӲXL�!xJ�»��9�c�������$��S)쯧�{��Sp;����@2�"�N�S+�/v�{>�#-�dO�y��!���|�߅��ϟn����Z��pC��2�
m ��۫��0VM����Җ��`ߐ��p��P�X��ӨDd��ބ���i_�1��A��#	��3����Ouu����~b�h���� IO�`ײ���������L`�cj���#V��vB}k�����"c�ޓ�OY����y���F9��e�(tѹ��fJ8����?��o�p+����XGh�)&���������X�tnk��R2"������̼�ϫؙVXǈkg���>�w^�\3�7�`&����Զ��Po����
V<%R6�0���Yn�]�0�MU��-�S~5���E�jgb��ۇ���c-�'��VV���	��i�����L�|֕>�	�b90D-�)��C����<�����B'%����؛�(�ڳ%�����V��U"��9.?O,��c-������}�6����k�9�d����`�M2��0�����A@$$5��q�^�C}�hY�C)��Y��AOa��X�1y@Q���1��x0,F/%��s�G?����� �c��ff9�mb�&��o������9z�"�����}'�0RS�� 9 �>�*�z��'�NrO�#��kN�U����>4�οd�9#�d�#�f��w
�-)k��}���u�ڙʹF�qj[�r*	����-6�˪�	\����洷/�bF;��|���4MNE��V�_����/~��p^V�b��˹�9�ʰ�Nn�-=q������ڼ
?�(��?�5들҂�)%��p�!��M!��+��YF��7���!�\ƣ��yY¥�� ��,����t�b�wn�C���ŗ�|X8Q#�W�c�q#@�Tʲ]��i�r�A��7�q��he�&�����a6>p"�+��_���U\�����oW��*�/�­�ۑ��;�J� ���v�h���m]Z��w��ۡ5ة�&�4_s��V�%�p������ �ƙ� Z��ѐD�)������i�>q���|s���z\�?${�'cd��@U����)^wT�"�DK,L�wX�C0E��	���1T5h��o=�6/�]����J�����*cw����^��(Jr�q��r��whh<�9��+��?�V�M�Z5������m��\m\����޾���p��͡�2�mi�8���e�_�B�e����쇚��u-xp���\	�2gp���W|�`�wOu�U]Q�a ��f�m��\���W�+��� �� bCB��[�y�;��RG�<y�H{�ƒ^HqoV(�Xс���WtsX(C�lkg�,��;T�aP�j�5*�������_�v���64�)��� �c�8������� ���wm& Z����� ��:o�9�{dcpN�ON^�?���L�v�:�ױF�E,�m�ǯ׹�KT%VS��a�+��y�VfR�S�ɀ,�+f�?e�N�gJ��4�W+��`{o6	�cG�3��}9����~�����VC �LS��^r~�� k��ڜpO� ����տ٦2����2��0���ln����v���)1��X�;POp�g�N����f�����%Xi�;�;:���,>�����]U{Ë��ʶ6�����a�����x��݉L�{�(��tC����Ƹ���D��1���v��Ԕ.U�����E�iڎ~Z����L�&��h�G���"��BNp�C������:�\݄��z��\3��M5k��\G��f_��������]�I��YN2(��@��'=�ϡ55�Z����b�XG��b���E�^�D�
<ɨ�֖��c�C�0��~!
���sI��aЫ����X;�9��	-�B}P��R�)���VQ�����v�_���z>�R��p��z� !q|�G��o�M5fD��.0��Q�8�q˵)^,�J:2B��>�B3
���]1~9��J���_����@//^�롟V�,�w��g���I'�,�Ҋ�Ob�� &�,�T&�3f�O��S�u��*9c*���Mi�MF�qK�w�< k6�@�!c���4華䈬�[����ZMI���f^>`k؞:z���Y3���Ӳ�' u����p��[�9"<(���z�����0�*��W�h92�%2���	`|ma�;�=p�[A�M�񎬑�0j��7�R@Fr1v8�pK�E�I�����d,E�	��ypͿy9i��)^Ļ�Fh��������6��j�5���{�F�7��w�@Z��$�Tc�g�/�L	������Œ��ʛ��8r��/$-��>��ƎE�Z.�r�~;��H�黓 }TR�9���b��Q���S�H�ߟ1\������������ҷ��*95D�n47�$2��ё+5�%�0��C����Z�e��/>\��nYx�yc�H?�4�"�e��%��<�M~���V�\����a�����1]%����e�����x�7;�A�5���=��S�2���ŀG���1 $�9[�J�k����O�K�/�!1/!�OW_k|ѡ�j����2�?#��m�!u<G��kAtb"���tJ����F�:&Qݘ"{�oik�`a�����'�$�$9�A���n�!%{%�¡�����-��/�y;i櫞���]w��d���տf���I*�Ԡ5�<u�8�7����Kx�2@���,���՗B%��H��2�����F����(�D]��ͨ�i"�=C������p���Mt�Hؾ�	u_�j�e��w�,��e����l_[�|��PWj�b���,�9X���f+��oII�2��&x=6 *k�y�6ֻ�X\^d�]��`�<�/�W�z����B&44���La=�*��h�l$b��9��A����*4(b���<a�!����#����=MJ��~�d��rYUr�����i��&j�]
l?�!2�.��L��ه�q���R�5���8���gwk�Z�=r�Tf���jM�=%���Y9PV��\��9fa��ȫ! ��Wt� ������ih�����[Zd���Q3�ɇ)	Nwh��M���2�`N�U�:ۖ�����:g��x��BB��yb7�.��9p��S����#6	J�ɿ`l�{"��pPΧqK�l��l�V��(Ʊޜ�R��\����l(���+d-ᘇ��6k�Z���^+@�)�!P�/�Tgͼ�h4��1ɇ8�����e!�YZVw��y��K8F��I1TE�w�=l̋���VQ�o�_u-��7��̶�;ۃ�[{9��U~�-ӌ� ز�h�'S�=f����xg������e��/ŋ�������䟚�솳�dx)��˓):��6Y��)jr��_��2^���m�ٷO�zh�VR�����;�����F�]�̣�q����oU^�YI �421��Ʉh� *��g8��K{�BX(���$J�^����\�_�AJ=0v��ɟ���${���-*�x�<�e��Ч�N��T�Q" 4���#�����n�T�����`�f�G��|Q˲@��^�������qp{F(F"]���M�����z�R7sM���Ĩ�ڦ�����pv_�?����.���pk/��C��$u��%�{d�7<L��=(��Q�/�G�<��c�V�y{�@z)R�����P=D��)��ȍ��YF��k�OD �p�x�R�J>SݻJ���v(�Im��L·�F�]*;���~v冥y;._�7�<��������=wU�5Y#]�_Tȩ;3��T�۹I�;� c߬�/��>i#�4��-�(�2�9)[G{~��`Uנۙ�p���2��ܡ:'��/��~��t��X����7��F��'�&b�P�!�b��ă�*����%�	.]Չ�u�O��~i�24�3\*����B��W7�B�I�����N��I�#J_�J�7з�H�Q�P�����c�Zhvx�n[���'˷�qO_�w
�ČATLu ��*��I�y��y�����6�Q)9�J`UD��G�s�\��f�#��z�D�i�S��ڰ�H?�Pj�{��(Y,I�ӊwC#��o��h{s!����ϦN�8`�� �o�B#����i����[������?�nH�yl� �(���Ӯĭk�|�C��x)�Ô�2��<t��n�XZ�W�u(H��>�S<� ����� 
�5��)N'��3l7Wt
q��a��|�Y��t����a���v5���۟Sٱw������IKG�IՎ���>į �Ph�� �(,R��3��C`Yq���ܻ_G����?Rh��s���^.���%��q3��炧Z�9U��Rk�M?X%W�DE���U�8�B\�Y�&(�m��.i[��/�&��D������ٻq�� |l�3��VK�6�u~�h廇@#�W;?��*\�c{���i�~��i6�_�� ��WZ7P���f�γ����x6���X��h���܄t��u��RQ@dH�U�������ilu�ޑ,Զ������8K�F����;J��ʫ��ҽ����!,��C������� �H��T�^C���t�ͤ�P]��2J�������v�Ω%`���e[r�*}���6�ΧW#M���;�?rx��G>���N�z�pKM�pړ6֕"�)�G!�� .�j/p܏��� ��y��oyAB�P�#�;j@�1c�=�7S�\�9�OY�׵��׬H�]s-_�?usiQ��9+�B⏓�c
�^kD�{��\�mV�ܿo��gx�	}�$�3����:��Q���$��$wr�bz:��c߽n�$�/�6��Rʿ�"l�?�����x���9>��Y/*[�#���_�И�+������w�Q�k:�@|��n{g.?���TJm��
��6�¨�.� )O&f;7(�*>1#E�7�T�~,͗�% @�]P���_��}�t5���76t���5����0	�~?��0���,M�s% �n��m���e���ܝf&K}ߟ�=�ɢCի�ɞ�R�ưF����杂1L�o���e�in��s��g��R�Ά�N�&� = e�geR�P�0�.��pOje�e��͆v�	6��t��'*��t�D`
ue]�̪������������'���r�ν�KV�%��̱� ۗI��u�O���$蹻L�m�wY)����xi�h��nѩ\��� ~[s���V&���Iv�"�p�i�uI~�v-��"�WYV5�<D�WCÝ�hҍv6�Y�j<�B$#���d �J}5�D �PE��!~�;�6�h���sg���ł��C���]�T%/��H�*^�Zn9ڢ��gBM����'���
t�IL9��pX,{|c.�PL�)�h�:��/����F[��3Ȃ������q�N��M�Ƀ�6�JyVq���o<�/���#��*�[�BF�?�����%%F@��Q ӂ@+��ߦ��M�W��Y;U���[�<RE���ks�N�
��Q����4<H�,�_��?�m�����9����3�r��7�%Z�� ��-��)�(�~���}�B��iQ�a��=���H�Xʅ�ֈ���D�#w�!������c=�٨#�'�l&�f�D�D%X�Q��т	� �/>�x)���C�c]��3�H��@�����Yi)8)�)2J���<KM�#��4��
�C�Ȕ���:[i�|L��ѓ\�|�9�1B
�~Jah �l�����GsR�F�h�4p�r�D�3���hA�r����ߧ�"�=?���'�FWիd��� H/�X��9��_�~p�
�k�Z�G��,4=�!A�����ߪc����Mn��<�����!\��w�(��HR$���r7�J���%l_󝡔��
�z��xv����//?�j�Z�!|�&s�%@����b����K�́���N��=³���X1���SEuv�ŷx��o(���D"�ʶM�	�_��=�wy�DS_� ���a�&���=}[ZSa_��#T`��&y�'��Sk���c�����������ͻhJ���D���6��;9W��O:����?��|��v�z�����c��1x��l�>m�ji���g��ڇ$~i}FJ20�n�2��XC�[?'k��|L�q�u�*�C��#����gX����eΐ�Y��� d-��&����b���z��>Jc1D���CXn38;U �rf r���PR��)�G��e��T�o�j]T���q�� ]Xj�"O�B�.�xF?u�!��p�:~�?$�72���W�y�v��? �*?�o�b��dAMVR8|'�Z0��uoN
q�[.š\���P��W��`��eޞ1|al�<H��>%k�s��#,tZ�1����#b^�'F�?��F���P�W��|� ��e�b>N-��j����P�y֦�B3���_���*k�-�_�9�o�b���ͶY9�[V��&'N����]�H3�� ;AuU<��nJg�4�ϧ\�B�U�z�`ۏ��bÁ�C�,
�jx30�#C*�2ZBa+���)�+$�պ��q�|��3s�����y��"D�4�S��kZ��~���F/c@�wJjb]b�U`,��j)����g�t撥�1!�E$����ڝ���(f�v��S��Y1�82�i�(��=�N]x�U���D�lM��mn���i6G�������b�u��M�У��$��lAi��e������C>�2�|$��N�`�9���b�Xٱb�\��4�^~t�����joq5�/Z�g0O�v�m&��!�	��Y�2��	�����~n�{�<�kP���-�h�H�ox��޺Rg`���������'����K
��y TJڤ�c�\`ū��Zӊ��US��t�9��B�5���rݤZ���x%	�m�)%2��AT`�
N魝t�X=&�2��K���}���G�G�_=�[I�r�ң�6upN��V4��:��7v���{�E���/eE�E}<�赌~�����P,߭��:��%;�SdH�#Ҝ�Z�?�{M�z�	Rs}�4�E�t��>y�3=��zr�|P�uT	z�r7���)@��>��F��&��
̺��;D���d;@?k>d+nr�OGާ2N	���T�ZB��r�U�x�#����}�V�/�<ʯX�3y0����BĖz�3[���9��Xw��Cލ8��E�@�_���률��Ҙ�Ǵ��4w�VdݧGC]�d���u)Qy�	����9��qf�sG~\�$C����>w=�^+M���bf=���a�As'��v�kC.��m'WK�>���Z���Z|�<��W��z��+�E��>�� BV^�V�A4�:ˀ"3r�|����� ��+�Ϙ���L��!�Y.C�Sq�v����X�g�>�oc%n�:�l&��M�FOG�2�*F��Z��G-7 ��C�^�`���DE��0�Y�0*dޙ��h�m8�q��ꚦ5�"����Umh >>�����:7��!�C��Ѳ�z�HImy%�HaX��  i"Zl��4�h��ͨ�˫e������~ι�E�K٥W���n���Q!��ɍn:�i>��E��~u��ǐ�<�mB��G�`M�5@�s���Ò��1�A
��x��2���ʩ��A�ɐ�B�V�n�~ %Ѐ?�-���U��uk -M=2߷G7��jQq�h�,���6*DG$�+G	=�\��F��Nw��/�Ě� t(�K����\h�!��sU~�0�v�����x�i�׋�݂�I�3�j�.��&c.�"��[���NC��\+p���^�lE�v�:��O�)a��p��/_�_��~m�E�̺��
5ܯ`
NG) Ѧ��a ���7��ه��\e�K(���pj��sE��s�^+�8���|h|�?q�f\�a�&u,���A� ,\�,(�p����F��gJ�o3"4񐳿g<AfF玎]O���> ti�)�,����Λ�q���#ó=�|ۮy���=�`�� �����=R3��ٿ4��W�l$7�����7c���Dp�H	B�%��|����:�ڢv16F-��i��u������{/�X6VGƿ�b�J�-��lH��Ha�����M�qZbT���!7���F ����0�9�+�Ϻ	���QC�O�����p������'c���t�f�1b	�i��	?���=�4��F��'0�^�\~G%,�?��m�P����������xI�� ����E+�	;��j� Tʖ=�u�f�i��y�'^�v�g�����kO:w�A�ˌ#���$����5w��.WT� a	YV��]d���]��Rs�i�m߅<���۽�.,�f��p�=zXF�j�An�S�R��\��LƑ"�Ct�/)����v���>'��y'RU��ǻ�������%���|�-a����dd�Q���g���%9&����2��ktA��s������2c��3x�8���lNI6��w*���Ȕ�0�eF�1àƓ����� ���Z�~���.���<{.����8.	����dF�����~^�h����ѹ��G�+�Z��~|����!*�j�c�'�q(�ru��80���9�&AW�P���z q{R+���7,�{��t��Qd-�p���'tJ�����p�_�ȂTxS���!�aPq�`����E4ŷ§mi~7v���1�����#o\04���]����V�aҾ7bKp7���˘�Le���D�J�}w
;W:��%��4�5��t�����@$�M�AwUDH=' =� ����]O��p<]]ZR�SH���Ќ(�͍Q�:�vO�_47S�߽���ҡ?ճ�̦߸!v���s,���+�$9�`,����Y&.��]ϙ�Kn�|�	�H��`F���z �TE#4�a�����(s��\�X�ȇ��b��;>
G����n���Y_�/�J�����6i,0KoA��{0)�WWjd�ft5�����v�U���?6D���~�h�~�Ej���8��V�(���ݣl_ �ɯ�~�*kU�"�W�_�n /�6�B�tD�KTV�:�}[<�rfT��;G����nl�`��],R�v�Q6ܤă�]Ũ0�46�ޖ�"�Z��]�ˋ��P��U ��(�y�@�]Z�0z���׿z�*t��s����F����Y�B#���}W��n�QM�-�U5D(�E@Ae��k)�op?�%�F)���V0<��}��� l_M@y�A�8[ L����� ">���)%���W��Q�M�S���>�>W� P/M>@���ļ�F��$��{�c������`��`��O��8QS)ﻍ�s�<�}:��늆���`��_ X��R�ʷH�I��T9�X�I�Y+�~���}
�W�̈�]l���_Y0��	4;�Ҹ`�,A�4��h�{�x�5:�aQX4W�Fsk�@ ܦ)�$	L�4��H���E�Mw������A$��,�+�t[d��㝗I��0���;�����d��޼L���S��A�( �8l]C힋��Ϣ	S�<O����W1�0r�����0�墬��Bx����'vYz'�M��ȑ�� �M����p��R�f'��d*��U$ J���~�34%{������q�N�� J��a��џ��@'9��'��V"�7-l�����Z=���	Z�y�L+��%B�Lk��{���2&��ɱ̯#�K
�r�
!cT�g��l��9,?��r�� s�Z�Z 9j?�Ǜ��6�x�2�4K�{Nh�!L�\Hұ��OFd�/H j��&$Z�Y:���D�.�AtYP�WR��O�+�!�E:Ⲟ�O�'���z;�\�s�Җ|�`��k.����,<�i�F!����X34&��\ �&h!�r�h�o홺u��`��H�bl�����z]���r��X�5����Po�����۞�b�����T�]�_��l�z���"$o�òWx�
�5���`�=�Q��\������E�WJ�z�����;�2�V��fa2d�+n���~|��{{7�<g�Y7� N��>q�E�`�9~*�����'�`�),Vg����cgض���YxxC�+I�O��N����!̇ON_��3`K�QG�&���3g����4�~8�J*{"3�hkx�U�BO���Z�Nq�۩�p%U=��dD������R͂gM�̔�Eۓ.��'�}eQ�{�S�S$"̛Q�3���*j�.�"���T����v��a��ȡ���;��9����h���Fg�.��
d	�Jx�X�A+Sg��@�"	@��ۨ�ǣ��
�P��7�_����C����$�4�BA������S��۹B%h��'�d.�V2��[�b�TLtG�^�͏j�����S�]%6��w�T���S��Gy�Ñ�aN&C��l|ȟ��o�{ACqy��{��S9naC���B��X��A�_����$���o���%S�삤|N����<�0ҹ��ý��I]B~o�>4@𽙈�df�rprO ���WD�j�v����o��!M2�Z�{.�o���BΥcMG���h�T�R� �0��8[�,�ǀ �p#����0����Qh�ML����r�әg7��Y��@��N��¯�?{�a����`����*!�%bK �����̓��6Pw�������BU� \�[��m���[����s9�AL@iS}�pV��5uج����<�И����V��)Q���M�3fŋA�������h�	�:�ـp�36f\����-�0�u��1�9k(�m�吝��i*-�����x��׶�*���L#�<�x뎎~��i D��Ts�a��P9�~�:��>��w�n�kg��f��g� R֟_�%���da�T%U]2(�!��rt�a�d�g>�����b�l:��\E �e2dR� ���W���v�P(͋���'!��#}���Jf��j����#]���B[5�.�U�A���},�ʉ\X��[^,
\~��M%|-��q�2힛�M~���V�N)���̶��҉f��!h�q��T�t�?vRhe��{v�^�GK�zc�8=��,���>��-q\ɯi����֯9#O�	��Gu��/���Xp┑6S}v"=W�4뮇ym�/oqA�^����ï�X{���7��/l�K��椐���{s��s�^������Y�Yz� ��4�j��`��>{�7�a���至���TJ��AՄo8�w� ���Zg*�[���y� �^ع���_���~͟�<��Ɉd�p�2`Y>	��9UՂ;�#6S��w2o�de��]tl�>R̌X�-��)�zp38��K��>�P0�~6���I�y?�#l���e�G��sɗgu�ֈ�yñ1�nU��6�9����� Z�׵�w.�zhչ�/���G�ܷ��y�]v�&7��i�ChD9'�W5A\z?">De8>��:> @�����4�jje>j��E:�;���܁�+�v��?S}+wJ}ʐΚ5�1���Δ0#����G僩���X�^��_�;ßO����޷q[�`����Y�04|���G��e���/J�$T�J�0�	xE0V�w����dD�Y��g�,14\�)��hgzX\��J���;� �p�G������Q=��ӽE�����by�9	�,ŁM�L�v}����9PU}u:�J4�?��~ԗ���o�w1�}�Mغ�Q��m��4�������6'5�oS}�/[�!a��Qu��\�*�������oh�W�J���h h�����K��l��>���î����r�Y��R�k��Y(픍��Zf�j$YɊm��$�I�%��!�u���f�(Ɩ@L���&�	'<�]��3:!�V�s%P���T�
�,=�>prS�0��>���s}_
�x�ٴ'�Ŷkî_�g����|����6���>S�<����V��̱ai�Ao�Gv��\z�ȵ�7��y/iY0��7h��C�G�`�Y���+�|�m�������T�njL��`�����v`?z�� ��`��ǃNjL��b*ĺFIB2" đ))$(S�A*T(�`
��N
�����Ō#ڞOj�o��![��@��]1Ne��.�utv��X�3�W��Sq���
��>#��oL����9HH�nf@P�!&��9RrYeB[epឱ�ׅ��}�X��i��/��@��f�̐�x)
.=7D
A�2�	:�V�e�o���"�b�����j�B�d?!	m�nX�$r^+c�*��Μ��C�6l��ɥ_����-�S��w��Dz>}��\�뾼*��X��L�O*���I�rje�`m�����ʡ��}dy�U�#몗�A�˫�a`�q�����!���ls[ّ!^'�~N�F
dcR_u��$Kѫ��RN1����G�/"R9X1�\^�!��I��db�+��&�3 4���q�~����5��M飞ʥ����J��'�_��m��U��=\��k�K�ȹ�qF�[4�yS��zU��k����2Z����]*E �~+9�&P\�h�)j��C�y��]ys|���0�xϯ��g\��O�"�}PP6\����y��W�x��?9�����_ᩖ�0���iw�fl>���b��h�La/APU�ج��Uế��	�o\z@X?Et�Q���ў��3+;���rv������2/��Z���g��}�M;3�$�*ĕ�U7�����t��x��}���n�Y���&+�2���u��$ ����\z�P�ᩊ_����$��շ.�m6�;�R��ڂ_3Ƕ�B4�u��{��cu�w��M����ޔ��?�/��SUA�̱���W ��<��<��S��(���f�c�Ž��;^kR�z��������2���.��"����Z�9B�̸�.⻚�vC������ �(��jUA���������:�u"����"��7�\�Ҥ!Qm	c�� ��+��1z�n���s��λFҾ����e��~4�2�h�c�R�d��M��_�c,�C��9��L��y㽛GQV���}�Q*ɉ�;��s�p��P�Z��������x�nu��N�B���KHܝ�Kj��*��y��8�{����?�<̗��2Џ\z�9N�/PMhN>��(����.k$e5�;V� �g�!9�.�,��$���NtM��Æ۫�@����g��U_/;;�P��7�I�c<�%�fj,2��g�瞍�M��@�s�'��g�Db%�p�6�v"e��a@!�"[���Ÿ�R���J2@�$ӌ�Tc�c ���[�1�	�_a6�}7�VG0-�v5e?(t0��tu$�à"���7G��ӎ�K�N\�� άw/��jcZe�aK��$���O��)o촂�^#���|�Z�P �a���/�~·6�w)H�U^ɬ��Qǎ�g&� �r[e��U��\�\�[�?},��.P>���܉�����b�ǃ���G��!]*Q:���>�,�Մ8<���c�����R	*�V]���3��uե����Y��n<@fxCJ��,�k4�2�-��=̾�4PǞ��֟kGi��8�`�˹��95hG�1!N��� �H��ʑt�F�V&ȇV+�`P4qy��E<�/�9��"�Dk����G�=q
שs!C�^�x$�MI^�Q���y�9����#*���"�fN
�˾�@��aT��]�l��L/P�n *�c�q��+>�� U�|n�1�٦ T����8טvq4�DN~�BӨ�T4���ߛ���`����	���!Ȇ�����d,��Lh��ժ @/x���K8�{��]�,�?:X�B����6w7�
�L�u��P3^���ׇ����R�&��\k/\�ܹoK����#��E�5�`�)�p�誉@����w2�WK<~�u�I�@�ӹ�P�4�g�����{Vr��m���Z���9h����G�q�h�f>gN�\��d��6���#�Ö�8������3+�5���V�%ʻ~��hpk�ku��g|';o���M�����EG�LI�p����pX�Cn�ȓ?�
�a\z)�v1	�� �~�;4m��d�c�D��p�Z.������:�at�\�ԅ{�FCl��X��l**o�O=V����q32O]GpQ3Odf�.��D^6#	���&����Ne)�@9z�(#g�m '.0�iOs/a��e4��<BC�df�k�۴�^Y�a����a�J�Zs� �{Gi�㝷��[A\�1f�Y�j�r�7!T�_�R�gt��;�=j��En
�wY��J�i:Qy�<��^7ˡ�ĩ%*��{�߳�� �� !?5�ƨ��)�/
���X��25 9��"�:�E0(�#�J�K
��OC���|��_e�SD�o7���#�Eϗ��m0��Z�L-Α�]���3��T����5��0��������t^yFC\�h�:�ņ�ޯ�J�kYF��8@����.�:�T�(����$��\�9�@���0="}F <I7�F�˨)���NVa=�v~�x��(�a��=��+	�/��*��O�;k� f~G�A�,l:�&��IA�{����ͯ��U��Ыorc�1C)䲆�����&9���&G�t
d���tX��r*��:�<�hS���=�Zɶ�Uދ�5z�t����nPx��l���a���qT&䦅�G�Ž����w��vUq>�����NEU�ã�M�\ze~�i��K�-S<�P�Y�xL0��^z���N�e�fgdu�L��)���䴗dXM��I�?�w������˼4jQ�ҳ��G2�u6&¥����?
�u:����w	ܥ�K��s�(�dR�wN߰D#�-�>�U��~ó��!��/�|�,X�o�L�eT�M�-<�C��>8<������$܂�kpw<Hp'���n_���s�����Uݵ��޵�)�DOJ���Mu{�, Tٱ�,b���'��*����/�����H"��)%��tZ�5r�� �F`�Ǻݞq��4yL@r���e�չKP#Cp~��I�g5;��@��F���x�~4�-~?��;
�8HYXM�^�r�K��]r�G$�Bo$h`��̖�!����\����e�k�=�%8��;�����u�OK�C壯l�;Ip]gg߂r�����jc�.ƽ��֛�#���o��7X,t3�P	w����|B0 ���|$d��u�m��D"�?�w��B���T�A2�z��q�`TQ�v[$äl���dYLt�B���H�EX�H���>�y-�Hx������p�)���7?��瑰W|��S�S�{��چ�(jO�ABچ>������˽��?��=x��E��(C������&���F�Ƈ�jB��'��v���x�p�l��hKu ����"y�! {�.3ɏ��xϙ~�1��X�09_\�-A��t9ѭݾ��W��w
��7�񥬶47��fM_�79N聁$ ���aMSº�������Q�~��Y81wk�D�M�uR��ܗ�e��Ŝ>=Z�I�����=�/�����G\N*��evs4�c�??�i:�q�b�+�� �ݺ",2�a "�#�VK|)R��%�/D��	L��9�]ޑD��?rP��Je�q&�ܺ���L(�m���xśG��8,�$=A��T�7C��#Oh����wͅ�g-�<U�(��Xh��Ɣb�����{��������v��M���u�a>�jEب��p�*7׶y�g+��'=Mfz�_�Կ@�hSN�Z���Zj�D���Кe��uȃ,G������ތ�Vz`��p����*
�l�wJ�fE�`�ۉ�Eu{6�<�U|���AN���Tb��rR/"&(1r�J$�ǈ�H�I_��sw�KLi��?s۠w=sc!
�
�EŃV=ʠ�&?~u�e����`P�\�.\��F f� d���Oߵ�HL�u�Q�b����qINAؗ#�d�h��0u����~��\�t�E�XF�ο��c��z�W��4�����ɟ���l���n.�ribP�e�+_{����q45ya;�΃30d�M���U���\���#<l>�Wf�UL�L8��iC�����ߦ���+�?�#x;<a>J�V����/PA�l#1͒��R�ܼ���`��;h��'�c��x-z�"JQ>
m�i8:�rE�X�D[�R/ǟ U��H��.��1��_�O�c��_8.��ٓ� �3��j�_Xb��I�@��=�Ҙ�9g���a��'fV�/�W�I����� \x�M�Ċ�|�%�2�����+�>�w�{���u��Gx�������2���B�(�� 2������D�P�hԑ[N�l�����h���%N�',��mY�|�նY��{�Y��&R.�n�'{�~�:,ʊH���cP�.i״�eh���j�L7[�M�B� oA�nnH���_Ok��hI7���X���bN����oj I����E3K{*�|�+��x�{�����׊z��iU���ֈj$#��`�>D�}����i�dv �P.ǳ��GK�i�"�q�i:Ht8��$��_m�ZH��d�oв�����"�~��4�f�s+@��&!?#�������0&	jD�*�p��+��dS'w�]^�%0uF��y���^��A�Wl�I�`|l��%p�	8�a�Oa����6��4�����&'T�]��a���i�7U�8ȊnGO9s.����i᮱��j%짶�Q�J�؍�"	O(�ʬ����m$���F"��f]N$����\-5&��,C}�w����zy?�|�KȒT�F���v�N��"�=OJ�%��L�/�ޝW� R���
 B�k���bf*;����g�c����#�>�������Ffk)�џ������Z�+��fa��O�l>��	�>�������阥8��g�l�Vʹ�딓��k��
���-u�dЀ���1��wn�����-=d++��{*Y�[�Z1S�l{d<�ӏ�+M'��?�J��!����W~����ގ�Ŷ0��`��g�vI2EN.� �!���ML���hM�1Ð�&"����u�����;r���G80i$�b��M��X�������vJ��_/Ƅ���il������Bo�[(�C~�э;j�A� PW.|����Ux��аrJ�.���%��g7�T)���W�<�?�#	ڽ�� ����l�����l��l���5g~���x2����D�ȁb�&1"<3X�Q���k��/J�(!e�9�?���˴N7pxfZ�>k�v�)UD١��q�v�I�e���8�N���lk}*L�(ok���8�����``��l�$����wi�􆎋FH�JD^�\�1�Jl�����8V����{����fS�'S!�F띡��w�tF)�WU[�p��X\��L��z�XqA���=�w���Qc���{����q�W����e��E�d�ئ�����β+5��DG��>�u�:>�~a.��T��#�{��j������T-U.~^ �])�ea�W"����p����g����<-�KM:��ӿ`S
�S�+��I��@�5w:��xcwYW�2Q*v�̕.K�hQ.~"�~��F��A�-�8gS���+���ت��or��m<��q������U4�}%j>�������/<�o�k�D��o�fm.�Q��y��&�F4��Ur���4�?0�|A��1-��	��f�P�(}�v>K`�Q>�|}�90}}^W���԰�ħ�6:� M�i�ߖ�\���o��L���1Ŭ�ق�i\���5JwV�+(�3LM�|��NL�e����`�K��n,ޗ�^�;�Ȋ�үr�l�7�����Y�*I� �'�N����c˪�&Cw�����	��EC%>)��F��,]
�7���;�
Aٞ8������=V����<oM��^��mKw�T*�{uS�Ϥ��+ޖ;O��T�i�Sy�3�%��'ϴVA�o��"7��=�o�S}�w���֥j`�F{��+�/5���S]ܩ�h�����N���A
���ؼ�A��W�K��jh�M�_Θ�$�w$w�j^X�ٴ�*)k��;�z`F�(�$�	���������1�`��R��`c���0UeK�ϗ$�V��)�􏻙)<�V�_�bB$���nڟ�3�\gk{u��+�)b0`�]V �ks����g�GO��pq�Wi�0S�@E�W<Kpw['�qq�>���ǔ��0�����ᦾ�*�����z�ս�:�H�R�qe�4P�_|h�=�v�a�u�4O���������0����-�0z����kf��4�V�4�TZxm��H�e�`B����i1 �?ψ �c�WT8="�%��a��Q*�|��n:�Xϐ�QE�t�D�%�F(�I�d�b=�=q��e�	9l�H���0��^�v���ŭ���"�8��Z��GwU����)��3�?�D� P�J��$8�"�݄�l)����9K��Q�O����B����ho!|z}�w!�{,����[�-�,^��*!]r��J�_�̮\��x׎.���n%ɳ��d�0�����UD1t���ղ�+�.����p#�M����*�ö	���US��vd;[ĝ��t52U�w�3���?t.o`���r�H�!�Sz���!�*Φ�h���p�fT�Söl*��|M�8B�{��Y��B��Ö��%�x�dgF�S�����$��@����Oi\/���݉+�Maï��S�CEM<������vע���&�����D��n����iMv[�M�V�`w-��눠\�Р_�0�h��u>:���I���?�3����?:���޾��5�ZΓ>���f+p6��&d���F��Q6َU��%�{H=�k�H�Rv"X����<�b����V�+U�(EX�xcU�0PyR~-->4�t����eb����H��ȋ�=7 0�D�r�k�&	G��J�d�YR�n�j�؛6>�9O˻7���x���m��~������������:ˁ��'�9�u��;�%?��o�5�����}#G=����,ⳮQ4Z�^�q��&R!1��K��JmJ���Z���l~!���a����t���tw�@��l���Ύ��-���X�g�`I|~l�^��#)�������v�p��i�e��΄6�:`4/c[�Cc.���3�ˢ�i��{{Q!J�}��X7[`�@�2����!I�2�})��LnS�ѭ���uس��nT��|����5~~��ښ�bT�퉔�=K.c��#Z̨ ��Jti�nba����w�6&���N�~����s _Q.���\@B*�a�V<���e	g�$2n�B��B�s=��p�!G����,#R��#���0-�7��W����|7��j�5�G����m"\��%�����&��'�{�v�c�<e�*}JN��]t�����z���ivA�g��ʖ���:��`�Hf>3�a�''�D��]*[��J�����"��|s���> Q��^�������m�������~Aȇ����߆���܁dw��yZ�ɑ5��l�3L�(cz` ;�ġ�ao&�l$�w[^��Bj+��i@/�j����j�s/}��Ed_9�C�ȍ'CV�)El>j+^�I_p����J�~^,���{��}�9{�j���u����ﯬ��q�`Óp�\�`�#�9�pRmdK�)o�C+)�dݸ�g)m�:��a�4.%��8����� EO��� Bt).����@Zcҕ�	JBc�����I6�-s�CR���W�=����A����09��P�k�8�qůK�s�]�a���Lw6���^�;��~q?2o5������i���GsG�aV���,�p��Vǩoz�&���ȃ�_���l�2:���7��HHHg4���Q Z�M>V`�C�n�nų��Z-ʢ(��t�	�t�}l~3�����6N���_\m�|�|�w�
^���O��:�]�_���[���=yH����8 ԗP�`r����,��J7F3���w���X���>�KO����Oׯ���F^��C 6�]��$����0D����@�,��c��5e�����~Aö�4�RZ�@�f�?��M{R����x���ͬ�HB�Ƙ~���{��a�͈A���)h�#�(F!�0�������g�t�ڋ��j��G�om��o��x���X���UG�>-C<,OO�B����5{�n��4��kܧM �(���70�ƤVq�d�.����fb�����4��6.Y�}�n� kޏa��Ŭ���İ��ڗq��[��o���:Tך�S;-r�'٩���Fyo�?p\���9�޺��;ϧ)����V�R՜&�1�ǚ���/s�Q��G5��6��7Y�S��&��LsM���iŤ�X�C*'RG+:=��Zol\�=@&� ��P��i��j��Kn�ӽKZ�$��>t��2��,1�<j�{,U#����Fy�Z��2�N�Y�)��}IӶ7�6��D%�����p�B7W�����d*�*Am�u-��s-��ʑ��_�?ύ�A��-����9#�v~w����(]$�*`AE�z�����0��UW\�O�o���i>F���k�":E���2���$��Zi�:���@2]?k�F�!\�_���A����p��g!���z�o�?�߭^�0����0�����o��wn�t���F"	�4�!��mpB����6���_��7�S����O��΁(@Q\�����u$*�ֳRߤ|^�b5�#�=�?.ny瀿������ִ�$�y��j<exW���-�V��6L�mA6k<آ% ���k��8/��D��p	SF����9��"�'��yh������&��Ƥ�;��`܇�f6�8S��e���K�SP"w�C0&��'����?Ð�W]�ow�56p�E.��s���S��8�p��e{|��7F�w"���د׫�8;��+�F��$5�	��Cs��+9lI�T�܅��ʹ�NM�}%F��{e]�86�Db����-A;�V�����Ba`-�N����㯓���T�|0[ ��ǉ{�˕oP���8�J���q�VD���ad����
l\o�������P�_}N��<3K����3���(��z�����;��Q��ܿ0�r�灾Ď���+-�4�pcȧ��q:�N�!��t�1S�����S��"���b=�/�w�Wmn�W�EQ3�d�����_UO����yP'�b���������`+I+<s�^����R���f�o?�Q��l��К��%���};�j���Y�:|����Fb�'U�����6Vy���=�j-(���P�����nE�\�T��vz��,�0�5!`��
���bّL�>���w���͆W�*�%���18T ����XS����B=�_'�:�Z�@o)Z�-�[o���5A�AA�A%�#dͿ��b��К�Ѯ(��)����M��2��r��[PH��{�Y/kF�F�+����
�� �J�L��K��*��N�ܮ�(��7?h�~�!��ћn�h9}�х<l��GՓ�l��̚����1����k��9�����=^P�^�H�t�Ǜ����+�5`���2�����|�HՃ��(����\�c�;�O�E�S�B�"�۔H�Kߋ�� X��͎L��K���J�/Z�ו�����eUۜ�mm�pmn�g$w�ڟ���}���i�(#j����K�1��s؜Ձ��	�a=����+ �`c��4�V�]SX7i�N�7��l�`�
�h�9���&|і5�2H!'����;�� �K�<Z?�OF�M>��rY#Og:�#��֥,������:��ٕ�I�i�]�G�s��Nd����W�pd��1�#8jm��2}&{����m���}H5v4���_]��� ��R��Ը�-��=��E�PthIg��֐5�6Z�y�Fi��oH�Ϥiq��x��^Җ!jm�ϸ�ثw�&P�7��BYmWr}�=���?rKs`"1�6�]�kN2�lH�0T2�p�:ew�k�D0�R1�Jp)0VBM!��-M��6�bܼ�\D"�ݮʏe>�����\QW\�p\��阩��?vr�39��fU���q���]%r����8��'�Kz�7F��o!� Њ���j�ْ��=��gzm�u/�-�9.���u�S
nmn���k;�j;[��'��喨Ⱥ'`��*�.�/���em��ɨ���R.l
ns*�����ȋ�Ż�ϴ!�t���:�m�e�E@H�������7��tRo(?��Ss�?�W4}��})p<>v��4Hќ:rr����!�͖�E"
��R�̂Q��Tú0��A�$�D���[�ӡ�'_�No�6\>���-�o̡�eef��wWpDR��
�wφ�� Q �S�#�@6��L�O�h6:�NՓCGR_����f��B��,��뺱��n�x31!.$����7��v�Y"��~�gkZ�.��_G^!��C��Q1%.�[θ��@J�K�q�1wԜr�t��@�gհ�cQ���e�,X:\,���JR���K."&F�G)C�[3��JU����FAt�|��x�/��j�"�=^�\]Lo&\$f��r'��[�Y�=$�􅚘��蒻6���6cQ�<�yQ�;���~�Ԥ$y�4t���O~�O��F��i5�z[�-d��Ez�����`Ǧ�fN*���`S��t6*x=�9|�<g,޻�7
h-�������.��\�>50���E�Z�d�{�DT-ɮ��zG�<�u�G|����'g�E̕[�ǟ�ӠH�d�7�;7F�?FuR�M/|�ኲ�݁,���펅��!�G!G��Q�������M+:�k��[LW�:�|�J�v'�,1�]2�r:�F7r�����cyfU�Ͳ$`3��1ۑ,<���e�Gv9)��C�_}��Px�k�o�vk����s~	�*y�H��'�ܳ�o����X��m�EYo���u��7^��0F!�O���'��DY��ơd�ֈ�<	��k��R��O�#i�;�ojG�To��kΥ?��N>����^ԭq��KT���t�
���_������1P���٪�ʰ����*OԌ]�6�?�v����!�kU�\�qo�^T���%&���ċ����$G����N��.pTi�-�9-���hv�GO�p]bi��;M���,�q�����l
l�ꀱ��+\!��ޟ��2����r\���[�0=��C|��c��z8D��-U	g��L�l Z�R�yf�k3C>�,�j�S.����\l��Ĭٗ-�N���#X4�>���ac�� �Ѿo�"a��%�U�~���Yɍ�(��g)\�#+j����&�>����j��~Q��J;�0�ᭉ�}o?�N�۷�tB!Oa��~��N�e4'+�6$�+�%��f�#qyG�Eęs�����),6g͹J�QVs+��5�����RH�i5w�Q�$\�s e��q������E�'�:����7�Ɵס�'�wR��o�����*o����d�+��x��vYf�*2��6�'0�\�J(�d &%2x��[���"��U���~5�4���" ��a�W�*b]+6G�	&I�~_$�D�HcN��!�1\����J����Kg1�#y���\X쒒��;����9.<z܊�SۄLn�ꝑh�߀���M��j1��ziq��lw�\[�ڥ�h�,6�t=e��`�}���e���������[�K0��6��Ǖ� $��qG �	H��]&��b����C���t�F��f�΢�W���N.��T�ox��'��GਁT9Q1!`�1�d𴍟}6RZFE�]�dU5{iZUc��Gj�VU_��s�Ե�k�3����y��7�\�A��ћ�}�8�I��T����J��.>�>����1Cc$��kóm�����VB��Ԓ˓��H�O��/rO��Wp;�Y'a�%�,��γ�n�N9������k2���ꋨ� �:)Z�'\��eًf�& ��M�='��<�^�m�����V�7L��G�&"�N��$ ;�����`ὤOëjI�6��i��QƇv�Ew�@^��ֺ�OΎ�g ߞF�3%�y�O��-���ά @:Q!��_]�﶐9�e�N�֞�so�ZKa"(����nt�w;J��#������ֱ/�B�V� ��w!�塔���J��ΡA�Rx�3�a��|czN�C6�X4�܈[�tC�T?�ğ���f��昃c�k��R����?O"n�f�%bd
�p�g�#�U��|�G�K��fڣ^dI}8��(����V�!���IN�!�-�
nI��7�@� 2'����s|׸������:G�����N�PE,��O~u*��=Z��1z:qN� @�^ ��(>�� �f�ȟ���T&� ~�302����{њLU���aR�]���o���o���>�"Z}|kC3�p,z��[s�����BY.k
Ƀ�6R_"sJ��9��&`��������uQR I���Y-�IO���(�rf�b=���߆�J}��6z�0��.�S�	�'��g������u�������X��5��-��M�æ8������_�!��g��̟U��e��_PU��b�y ��v�߿�C��us��nCm}��
�ƀt�\2�t�y�Q�Q��i9��l�Vŏ�ԝ���Ha��_���T�ac-t�U�!sE� ���P��yķq�8��LB�lf�5������,4�-��0Y8���0&HʟS����;�j*<d����ȁ֊N{^':C���g��%u4����Pl/�߼~ㄐmؾ�H�bNU؁�&W�0uqL���P$��x�����ȥr�6����d�n������w���<���DY�r=nAՑK�Tr�cx�������}�z������T �O����/�.tC 7���z�jZ�:/]1� �4I���BU]\�t�����]H`�˖ �}��������MxW��o/���������O��R5����3V�k$ �{�>*�������@�;�H�x�	� /��������֏0t�����Zw� "�X�(a1M�Q���2@��cʸ�e��W����r���䘫A��4�7'��u����ޕ?&+b�F�A7R�M&�A�Q�4���z��N����"��_�G��� Z�ar<��d�GՏ{��BXZ��%9����wP�JKɊ&Xͧ����-����c�D֭�ds�	@w� L�I.b���V�]9��1v�Sđ��d�-ω�M�1jy⁆�/_n���2C�
0!�	L�@B6y�G{���p�U��=���p��N����5D�:m�[��ܜlI���Ud���;ޛـ����fàz�d"��&�.&�mA���]�xA�bY�U���
A���e*:?h��R��3��Q�rp��"�NS���������d���z�/go�5Zᰄ���&k��NZ)��-A� (c�"7r��P��?{R�EĮ�չ��:�K�|m=�l'������hv���O�̦�6v�{)�(k�bl�D�f2A�����\�9��Q�/�%}��Н���7��+�;Ɉ�bλ���ƭ�Q�.]��d�2K�k���c�����?�.>�«�EjR�Wwϟ��OɎ�Se�~�`]=��[_'�R.V7�M�l�IcH��?�f`�L���� ���?�vG :Z�C��:�rqa�}gL�변����C�G34��w6�����J�z�I\�j��.��������[���&��3�עB�*����-�	����"��zW�;��5z�׽�ܰ��g�i�ьK�ov�\GEc�
ȧ�ݷNؐ��,�`��.܎ж�����L(U
9N s�L~F`��>�**�|���MYn����	�tTPc�@KY`;@r@%��d�BL������{��+��疅�'���'z���-�o�x���6�����_����Ia�B��C-I��9/jNˉפ�2)w���.CÉw�>%0�G�^���n����H�z��rG��5�R�Y��m򉶲2.2N�����O?���i�� ���b?��v�l<I"�U��a�xF�mZp@Ih�Ks���i������A�w�-��3������}v��KCc�
VE;Ͱl��<ŦF�ZA�٠�P1��C֗ϐ�`�P�W�x#ڌ�Z��W�A֑c+|�EL��K�Ȕw�o��yi�A�Ԡ�ē7���p�������䊲em��9sGR6IO��U��դ���%��4u�M�֨f�M�V:�T����cd��A�#��\b	��q:�
�e�Խ� ��O��{;��96�/�z��柝=��b�V�����Z��}��@��&<fZ�9�Q6�Љw�f6����~��?���OD݌6��D��%�_[��)xl{��B9��T}(Ej��A��w:a��fTe-�uqR�=8A�^��h��7";̶<���1[�y�kxX�W��yik$^'\M�ܪ-i����5���+Kf��:�[GY笠��~�k����'���\��"��QD!���#��'�����b�����g����q����H�0�0��{�T�W�lQ�Ƌ�=_���y�e�W�7f�ǯ�>��O8f��eSv~�[ZvD�dH!�
��\s8z[u/~˩.[��\y����u�����SR3�`rv�s��Uu�>��2{+L�I}5S=�&�!Ƒ����D��^ŭQ׫��w*�4�⡽Il𮗬���;�Yw�r-͟e�sbŔ�gm%�VU4��'��&��rέI��ov�P���O�U���Fd_A��G�I�f�����d��:a:5!	^Spna���n��~�R��$H�f���l�E�}FY���)�I�a��o�
������@�Fz��zz�Ǝ��_���3�����JgX��aV��3�f�?�Q�$o���E�{�h �G����qI�6QKU���@;�h�qPF��kʁ�j�!�3T�=�&h_YRȘ"�vӊKBU�3lG�n�N�����~Y��:�?������vI���fR��{Sɕd���p"�����Q��պ��O!ԍ�j��t�w���ː
����Hg��#{�tg�x�H�_u��"&؏�Ah��'V�����}y�<�G�e-T�f-n����{�\k�_�F�d��s��;���jR�������$'i6��O�U�� )��w�^0�U�[x�,C`D3mƕe��$\ҁ�-�LR�x��h^�'Y��W��.WJ�}d(�e�kr �6�G��|�Μ
9�c�.�b@�=r�&p C�*�c"�.6��𭯎�tH���֪{M�_�ೆ��g�1�!��f���J%J��`2��U�+c>A���;��Cmw!	 �J[l�6�� 3$^@��ሃ:�S<5s�nK�cN�4��6Xګ}��j���Ţ�����7Z��:F|w8�4���c�:"�"&���� $�)��0��Z}<ޯ�����ݔ�u/2b4�B�-��eM�!|�o��s�^���y�������0G�N������	�t��S�l��h�M{6��ĝW�,)K����+t�ɚ�B�x���9u�Yϼj�|;�*w��N�A*R��i�j�J�1�0i��=�d�	~��G��P�s,�����ys8�+%Q9%}6��~���^�BOZ�n	���`�ԋN��!8�U���!�0�x�r�,�,�q�:��hIc��o%
��o�Z����I���̙w�|�٪$�jw(�z�w ��yd����y7�=�����+j�騋E���W�cy��:�m�&T��.q���N���ٛ�ױu���9{���7��ދJ��Fg���Q������L��ʘl���ۑ�
6xK�e{�i�������� ({N���N���N�0? c�3L8-|rH��w�{E��e�+�q��@�ql6��)p��:���j��+�̃�2��y������ַ�4g�z]�t𘆃��&ꕨ��&ŕ=�Ro{�-�n`�� *f�W�j�ʊ�	#Em͠/<e4
;5�˾�H�^	�FW�+^-�ZrPxղf�g��2�a�0:����ϰ/P�*�4�Y���%���l}�U�f��MJCqѢ�f�������?�;�-��`���8���w{��{VN;��<��|��V��1�è 3hfs�"���1��<E,6�G_O�	&ݱ*�)�AֳE���c����Y��{`V�ŉ�]�C&g�u���z!k$M�j��n�J��8l��2'���x���۹��m�a-�j�.FO���*��<j7��x����H�n>ٱ�ȜC1`��!ݨ�v7W��_� �4�է�o�qOGk�i]��w�h��A!��|J�5����VԘ��r��ٟE"�"l���{R���C��`\:�?6)03���"%d�n�Z�C�5�9W\�|N*� �����vb���=�
/ѻ�Ã69C�q��u�~�\���] �MO��S"�p��=����A�&)2[&kpE����G��`�DQ��^���¦����)�|�)��?6�N=�)��[R^��:C�K1ť�q�{�9'e��S?r�3���>Uh��6N��z�d{"�0w5�(����`�X7�ԣl�������R�Nӌ�iQo�V�B0�,��u<Y�ԀDO_�rj�����]�>�7��I<`_�Ơ�Ab�[tzgB���*8N�J�h<�b���p���_3�ߧj_t��UrH&����#��M}jt�ِ��s�t}��������$��|��������䤈M|S�!�6��y	e��Ь���`�!����6����>�O�
Q:�5[B�nb5��+��Kf��|��j����j͠",��r_�;��B�S!V�����>z
,�\Tw� ���Ey���n^|r��
�q<�������Ϝ�o�.h@�lH�� X&�zW?����ṔD��h���m1g�)E��[Ĉ#��"�bW�U,H��9%�s�O�t�h���B���0�<'����مqU6�C��h ~?\2��}��AI�dDc��X�4-l
;�
�~4�myY><�ٹ�0�^=nVU2w�M��2)���N�rz�m���I�䡚N���W�ܼ�=H��ݹI��5�$7�0�m�PJj$_�J�y�t(�FkG�j/W���?��=�F9�%!C���\Y\�na��M�
 v��]@¨]�'}
��3%�f������hp��m2�ԥ�������Y�t����O(3U\��Cl�r>/Hy���� EOI�#�TU�lԲs�I�^|:����Lŀ�*�O��/�FU�|I��H_uD­,�ֲ�i�ў��]�7��Q�-�`�Oy�(����z�.O�%�I!���?��
���>��RHC��{�*�Ͽ	���sȿ�u�|-7�`'���)��ᚼ~_yo�~7޲/�q&����C"R�x�
0���� ��m��죿�/F�`�G�*�Q����z%dx/�7ѓ2Z�̋�m>j�Y�n#�W�X]&�����HF�w߰����s��DXĒ�C_LGc�`����_�O��B'=�`�k1�U��qV�&Y�9zT�l%G��a�A5��E;�_�av'c��h�A�)T�V�t+
��d�R��;
��~N�K�γ�������^x��h1 }G�9���aU7�H�i�ܝ/}�� ��F,���`���H�Y�	{����Hz��`s�4�>�<x$�޼�K"������9�#��ǅ7]�m���O@�g�;�q�a�*Qm���Pő' �[ݸ��lN�5�!�N"�:���3:���ť����%��I��L�+D2M��r���<~>H���$��@[6�qK(8\�}Д����8Ļ'ì�k���_�J��=�U/#$BE�L��-f*i?�]�~���n�S���6�y�q_-u�O
K�V�ϾC��o�NcXz}�b�>~��.3A��b����M����y=׏�Sj����ȉ5/��0G�ՠ�8���k���|��z%�x�����R�~�-������@eL�μ����\�?�x���E�E�4�?`ek�"��y!uz�*8d9'��gu��Y�mp9�̈��2��
 ��͉ʍQ6�Ư�����fu�̗Av̗Z�,����1+Մ������ 2��o��;usJW�2a}�� ��V6r��1�H�N�̔�ֵ�_wz6B^���?�	�uw.��p�ӣp��jc���m��	dVkI����� dDI_��`�z^��^ǨgGm����mǋ��+vVa ���Ao�<'��S8�(5����m�2-�|�{D��))9�����/Q)�I��1���J\��r����ST*jܩ�_�q�B�>�H��)����F�j��NDI$ރh�2�$�_ @Z5�<��E�*���Y�4E.�Qz�d`��28ӿ�B������	RY#�٤�`��qx#�#��K4 � q'�ٿB ��4��L�|_���ջ�J�W��d�+���qq��:F�8.$�L�s�2b�ǧxD.D�;*<1r2�\��}|X4}�{h1}�^�W���*����1vBh=�L��i'����Z�� �R�[[r>mL��{�q�ѓ͐���*� �nA4�}�=��h5�`E%�cB� �'x=EW8��3���k
*��7��h�\]$��D��g^�����B�I=���X�pPD]�'%/�*���Rn��w;�/��E#�o>ؿ�'���u4���0UՋw"����җ��+�d��?���n�L�Z��3�}7g�٧����a
�: u�u��v��@���g_�^ O^�yQ�b��΄-�B]7�".0y5셭�x�4C�8s�9�� d�	
��Sk��S�[�X��8��A�|{��+�� Z�,x�\,E�!�t���VI�-M�5gi�[�oc�*,!���Vd���5��S\�V�Z=�����J^�5��Zx�\��H�e1Z�r�3�z������.�����9��	>Vr���#W������FkeN�%ؼ3�B;C�[�� jT�G,���%D���
͚�;�Aỿ�[{x����i�E4��^{;\۔���Mݥ
�M�+/��ϢϛbE{�=�K�C�TE�+�0M���!�:���_/�3 ����Aqu��3@��A�0xp���� �`����!8AC�����޽��ίs~��k���}�kwq�U�윗�����}M��M��DEeѫ���y *������[l,�sW�����C=2�u��qUFй��X�9���O5�3ܻ�1N�[IR��+�����W�2��ug�n2�Ƹ4�M	ɂ�)��%4~�j }g|�|��_lp�E>3�!Hh�fm�l-��\\,U�;��5�I_�r9�De�κ�-�BY�����\�ʈ$�)r�有P�o�Ó��,,Ж�m�/��N�% �/
Yb�Bh�x%5:���ʲ�O���2F�|��v/�U�,b�ZS"��{�,���>h �o'�]Ll��q;VPJ�$�ǿ�g(�����Xm*��o|A�4��g/p��)�賀`F���x*c����0Cr1& \�3;~�J���if_�ṷ�Y_4�5�$t2�fޛI9{��	L�Z�X$0(�Q#��)���.�X)R�6$��IZ�V0`pZ�k�8�j�|���1���yf�������O�>�3� :�2\ށDr��rp�^ݭ4i�h`����Ă�9��d�ah1�D؏J,�+4{��pӃ�\�k�k� X�78'8=`-�ι�W=� 0��1�g*	�4*� 8�^��և�$��G�W��ْ+l�i3o��@v�����M}��s��ciz$��#�yL@k���{s���:��Ƞv��~~���kE0ޑAz~h��f������ �Â�z�.���jQ�qi�YS�(b�3�}IKN6�.n�x���DB�f�"G�*�O!���9���9#��m�IX`\{�Φ��[̆2UC��ޘ�Pzo����E��������g�)	�00�N�@|w�z'�é��i��Zw�w��l�h�TxNj��VO͛e���=�����^L�,=A 7�ީfk<2f�1��������~�j����M���-������/�C�9��|�{g)��\�&�3�#�)<S%4��
R!������a�sދ�'ƴ��.G�'ᩳ2ұ)���#��:�֡�  =*R��14�<�3���i�x"o�0�(h�����] ��Z[3��}�)�'�|;t�@ �1�|���z$�7�|��qZ�]�����e��x��[]m����|Q|�D��W� η��ҳ��F7fǞ��aw�7K�\U�[������}�FӴ\\�A!��ӰM����H���3�;�z� ��G'������p��-flR��X�Vܿ"	����+��M��5�$��EzWɮT�o�yГ󥱰��1ag�7�:�^	��y
V4q$0_(Ŝ9s��CQa�i5M��\����C�����N��8��<Y"�
;ٌk�S�������z����i�3"F�ȆCSa,pC����b���(������T���B��gj�ʘ=�Y���$,I����9+�-�����o�J�L����o'�cQ�1�+M�3�����Ƕ�`�*=�'�G�6���$�1-���}����=���L	=�8@z�e?���-i���L��&Ǆ�~�Hl�u�0(���-Tr8�@���.�;��	 ��:�NR�������x�R 1����{w����k�o�l���A=	�zH�0S�}G;� ��ؽTM	��@Iz4����pV�ɋ��\|H��l"6�9yg�`x�#KUۮ#,T�%�M�k��T�kXp�Q��ln�FC(�I�3�����M;�R����ygM�GȲ��w��Ӫ�������.�YSP�)@�ym!MvYًA���+�B4y�������j���P���g�W �p5��n�U��<�NU ��`p*�qe����QǑ�Ѭ�����;�kK8�0���NBgB�r�=S2�gWޭ�|�Մ�u��/�Q�H����t���O�d�n��,W�5����"y:��=3�cvڔ�x�}�6��A�`*��46�tעc �_�������1!���Q�Ot�Q)
��������P��\�x�M {%�*#��
�4U,}�=���B�T9�;�C��F>=�FG�q�~-�H�.�x���|8�q��+Q�2�a��Rh�n�1�Wft]����$��}	5I�YG;�b?v��f���j�mX�L��w&��c΍4�0�ѓ���.k��o}�IQ�<�`s���_�]�����`���uڈ�tfࠂ�}%IJ/��`zw����-e��j��&s
AW�`�0���� #\�B�Lj��;I�uH����[?��b�x?3>v�G���w�zP�Q����d�#P}𐘪H@�XKJ1��/�����	��Yn.��c�
`�N��$:�Ɉ>��H5��}ώ�x�s�S<?+�9m��DEw46�+�"�W��&��?GW�g�ѿ��wX�ڲ��2�$��M�������������oL�� ���=�P��Ճ�
˦3�w�o�e�P�I"֫��I���>�( A�5���n��&��/v��~�Gn'���M�u�5�U�☢��4�]�蝏������������Wnz�Y<�L�Gq��+m[��@�|wywрڣo"5R�z�m�׿�M����>��s�
�pHEq 4 <4q�+�{O~������`Z�����c�-��hh�T���k�3r�Z�8}�8�d1[[~��vӎ%�M��f�h�;˳���o
L��FY��Vo�Rs�"_��G&���1Rv��A2+��0���-i��@%�=�늋BHHͮ庛pq%��
fd.����/ǘ8�!�8�k��˹�E"`�"'�!;98	d���R��TJi��Bی�N�柸̑��j�[O�fP��ۅ�{���2�;�yne�	��KLK$�����RT�)�q�NH+W]vd��{�:x�2mv����2���Fr���_&L��be����/�"
t�;*P�ԉ}��P��9ۑ�
)��w��XQ�@ۦ%'��_��W�c���	 R��в�����-賺�Um�(� J��*���r�۔Z�2��j�Ԋ��K�Ϗzv@�՟W��V��]���Oo�"��e}��3�A>��U����\awy:���z�c�����K�8����Bl�i��q{]ԧ�CH���Bo}��s�Տy��9�Ti\��5�!�~�^�vBbA��k�5ΗE� 8M,g�
��5��n�$k�F`V[w�)>�+��A�����Ĥ�b����}���ծPXSe;���؃'$�$l����w"b	���z'���Ĕx`Q#��s�UO�a�[�:��&ز�{cL	c0�5�`'N8oB�N��=%V�"�Rvc���G=JO���m�t?���xgb����6o�}����@1l�y���+oz���&r�ݏ�E�vc�L�S6A�����l���:K�^�C�J�PtƅHҍn���v�d����Z}e��bd8s5��x�~��*�l�&w8@���
�B��We�f�K[~QֽGΔq��y.���Ǆ��e� LH�C.k��Q@ŻeV��w<vG���aDI�h�HA��'A§��%:i�ف��vO�q�d�s%�w1+�����r��.CE��dQ^X77�o�(t����|� !أj��"�I���-MR@P�t���"c�Z�g���+G����ܑMۥ�b��+)����uD��
 G９ؒ��ߵ�a��E8�<�",OJ?�h�w���F�������vv3�&U!_���Ƀ*Z�4�Ǹ!���Xm�,󣾒2=伕~�-�\:�[���3�>�`X�$��l�wkt�y�ݔ�~�8rG��c/8:�M�5������_�Nf�Z��%F�41�ߕ?*?I���>��		�%ԁ�/�}@`�^4�a{G�.�F�8ğ$zDx�@�5Fx�A�i��J���+0F�S,����v&�
�*��H��WnE�3u����k��f|3���z�E�u1��d{,U�_�6=p� �d�=aKH�-ŋ����<pnS��L���3+��n��O\���6}���dV+K�j�(���Ges��o�Aq:2���|o$%�./C�c��sC�U៩�[B%�i��w�K���L��ddxG`��
�*�1�3���A% J:s9��ط��s�q�����9�_��2#�c��0�g>p�`�Y����\ܬ�P����l[�m�5��_�VR�~���0�W�wi�m�߶��2H=�f������)�8.`xO�x�����I���㩴�ͱ��C����*�Qb�Q΍��T,xE��m��K���X<2V����0X�ui0�qV-�FE�"*�,*��u�;�}�}�s��`���ձ���Y�+d[0�sW�j�ñd����z�>��uqR���9���>�tGPx5���7�v���,��I1���pe���e��v��
N�V@�4G�>&z�'C����'��-�����Ȟ��_�9��ɜ7{F)��(���Y<6���3�Z�`��4R�	��y�9��y�<�� ���}(�a:RL4I�]�[�����"l����L������ [J�8�g�5��,c�,�cmd�6�(o�U�H~D�HǼP�E��#|4�]	U��{ ���H�/a�P��,�!����W[|�{E0FxS��R���y�}z��F��0�"��4�l����m��BHG���9�J�?P��E%�G��>P"��7��	�s;�N�x�`��K�.�!�W[���)��Ee��7_�����LP��F ��,F�KH�З9'�Z�v�|���ac �Sbcǜt�p>]� �\fK�Gx������{���*!~�˸$<�lЕ�����z��v��9>�e��^�hU��7��������R�p���o����D*ڈ͓$ꭎ�ܭ����{�<��F�l��\�/��e �F��-�(ӟ Au>�7������h�ΙL�齲�z����&y[P:a�`��
�Y˅'X���*��{eJ7QP�2�.R���O��N�߭VOY���l�G��C�	IMCS�=�]wT�pG��(�d�jhag�Z!j��t��9�@'`�+s��rwЭX� ?T� �
�Zr3���$:]m��k�ݵ���,���O��0��aB��A~���B�뛩��I�$����#QU��D�V� �	N��ҁ�d�
���9�f, �v�[����I5�	��t�/~=�a�ng��]�b�Q��x�����
'k��W��&��Mb@~XYմM��yl���E6;�k�X��Z*e�lp��)N�|�Hj}d��\�b��/b�L�v�|<P�]AP���1��-mO_��2��Ժ�3�I&s��F�g|&�{kg�@��?h��O�Y)
�'�J���4s��L}rgYh��?"�O��J�sy}�3�*6���R��F�v�0JTe�����Xg�q�y��[V?���X�s 5[�G�E�K�6�{�{�I��٢r�G�ϓ2� ���0lx��H�FM�8bg�_zjO{�[���\��1B�uE��_Y�=m:<?�\{��1�i%3L2<�S{4+��Kv� w�cG� �I�t������(`ڋ&�C�l?� ɑ�9�_�.���X��qK{L8��vh~xb�~��)��:�#�h����<&��;����pzr]N��ɻ���/���oRD�hF��]���F�%z�ԫ��mt~��5"vJ,Fx[���\��c����#'�a��I�R(�S�Eq�.�E6���@g!	M��Gw����s�UD�v�ZNZ���]��X���d%�cZ!Y4d��������!�fp�ƒ���칻L�Y�S�Q��b2O�i;���>Ǹ��8����3i#a�˷�G�^�wC���.�����x�\.��'@�#0��qȆ��#/X���M��o���r������v�Դ++E���E0��P�p}���'�̒$�eӳtC�p�N~\7��Rl`����ۡz�Hb�ߣ ��)|�ߕXk)M��{���<�/�+��I�=T-p"l&�Z$��vIc�4�_?�ç7��m��.-��p�� �ouT����eLcdL�l�q±���.8�r��;jW�#�?B��Z r�Ы'�k���Kn��%�0I�lq����V|�!�B�Ywi�M�h����
�i�P��Ζ��j}>�[��P��`�?�h��/mԚDq�n�hF�ݸ.‖Mt����v샲$(>�<`f���������ٚ�|g�~�b����C�y4�G�go�f��,�$�<�Fa�~>7��^��߮,�=���
oR!U	#�L㽩~���rHqT���{|�a��<���Q�?�
l�����Fx�j~�|q覄�Ս��a���\��Eq�~ :V���m�e��".n�rS�n�Bc�.�t�M
��M+ʟ4[��0��ow�3%zޖ��f��[e=r�A�Ăj\(�����W�ln��W�1�"q�n� @Ȕ�_\��e��m�(��cBqFcv�vM��"�'�|�"U��%[�ZZa��(�{$C��B���5�D][B�����ʄ资���;ZA��_V
�ϵ0���o�<�����>o��;��Q;��HW�J4�R��*x�z]�-�^���Q��T�.��X$"{� �`K����HD���A� P��:�3��]Ǡ���L����Y�`��O�E/�T}��GdIb����~� c)��*�{]�J�焄�`���d%��o�ovz���Ӆz���ڙ�"�MbJ���ԛ֎"���	��<�]D�2d`�:�2�KճK�',���w&n-%�fk�@�������a���B��/��3)���.�"m��s�pT�i=Ϊ��g���as���+�j&oA�}�{�Ѕ��������tu|�N�~�<���`�(?���.��Dw�i�7��WT��X�}�̗��Q�Uh:T2/�v����yR��ܣO�IO<�D���%�V	�|v�7wba'�{M�yg ]��3ԋ��("�۶v�m��.�uc=+�L+T9ۿv�}Ы�"U��N�f�+�ID��|'�KEhW�X�H�ch�����'�o�|��pM鎣�eR�Dm����ل�H��˶Bs�x��!���s=ӂH�K�q����`�N�]�ġl�h\K>�v�Ȫ��'F��C8�I�C�>������s++T�Լ�RS�ɭ,#I��n��ɚD,Q<���r�ۯ�W4*�j�%x�Bn�g!ytKO�M?r�z���ʈ�)c����>�dP/Ip�~bZ�1s'�؉�E`2�';(��I�R���[��o���Y��[H�:�JMu�~�ى�k��Z���=�ڋ��AE��/�����}�F�:�D/�1���Iy�!~������hH��b=Q�-; �P�mo}��ι(����&9r��6�K���Qo�a��2����^��f���p�2������g�T�l!#�u#��⺮��	1��W�%&��NH�\DSh|�_��J ��E�[;Q��4��g?zR�S�Hr��I���ͥ�`��Տ��1��W��c,u��fДz�U�y��Gxk)�4���f'ɿ�0��2c��uΒf��*�SP����s%`i���z�#h`��RWE�>٧}�iQT��_�����%�+��٣�6+�|m(&��bp���}u���?~�x��]<[�c��[��&����Z��R[)a��$4I�����V�L8{�,�A3��~-�I���Q���7}0F �]�&)V��._��F%�`,ErV�(�R���*�{�+����^YL͆DEa�p] ����b�A��;�@Z!��1Ak��r~6$$��W`
�r��:�&�3N.�A�B�W���nG�Ȇ��*(ZNĤ{��\11
�&��ܰh6=���?�n�O81
�G#	�]��z�C�&�L�d�f-�[���Dx����0��S5�����ϗ�(��Ή���K��v"�e���d�!
�7��;����`�.�Y×�.:�n*�r���2P]]ܿhh���Iu�#n*eM��E*��Y}μ6}�kl6����������vt-|��I�׃j�3®�
�:���_�Y���H���Lܮ�k��cy���+L-��t���e���CK�A ���mXQāb@^c&��LX�&���<�y2�I]�Ա`��~���
���(�o�qKwX�ؠ���٫E�)
_�38r�L�m:�G�сV;l*a�VF�u.��̾������������]�g㻇7o�}�&�q��%9�:~�y�����?�9C�|�� �����ľ�}��r� P��Q^�͑|�Z@nZ��#�������!fpQ�~�h�'��t�#\ C)`�@�j��i��o����Э�jA/��_�/��G?��W�[۸:Tt졔1�c��#iL-0�\�}��p3�H���g`���TI��*H
���n�DȜ$��0~�}�D���DBv(Mˇ8k}Q���df ��X��l�Ww+����_Jm��h0_��MkUԟ�ga�?}����@��Vk��i�<�.�C&���ဂ�'�E����Ec�tK�J�
~���	���>?���-En�����R���͂l�{!�Z��oZ�� c�t��� ,�ƈG��A�{C3�"4���޲B��D�m���w�,����LM������F�� ��0E�L�}W	ń3��Tj�g�����g�|b�gBn(�k���V��� �[�s��A�%�^���:�ϒ�N���cY��j�$��$H��庤�.��N��^�v�\���3D��tp�_"	lz.���������t�v�R�C.�#w�@���R|y˻�#�'b�͌~.����	]2�Ɇ��p��I��zw�#�m%֭ʵm��D/[@d��^���`�ӻ3�86�7���@6���C�(�4�-F�]�;�p3>����"k#�ݘ�܃�� s��	��t��$5��8��VX
Ϟ�x�bG�h�k�$����[��0�-밄lM*�������,���mV|�i��dC)'y���
Ot�xg�tc�u�h��̧�ժur,��͸`��G�����ً?fR5.ڕ/��
����Q��Tŋ��|V"׉cM����T����K]"k]�������a�l�l�/S��o�r��+��<p�:���bufJ�)���={g4*�����S�o5�N�}�������ek�d8���P��N.�9���z�]��҂����k*w�^i�Pz+}�e�D�mz�
˳��J����@;�R�z"�
��!r���". ��B:�����?���æ'm��v8I;�d�W��Փ��a��̉� p�_��=S���\u�3G�_�2�g{K/g��w���VKP'��T"1dY��>��&]�G� �O��f$%��9���/6'��������t�Bĺ�[3:m��_�-m���Hm��?:^w��/~ET@F���ۢ��	a�aH�-U/: �Xz3�ix�+�/��~z�-^�u�O�a$�ІZD3ӡ�YD�Dg��I!
�L�,����C�[},{����9Р�:����}t��?�E�s���:ȱ���/To�3^��qp��5��@ږ���(���<���X 0�����@_Mp7� UA ��x�E�g�������oh*��b����	Ԗ�5�D�1��&S��o���_��X\*ݼV�����͘p���g����fSZ���y���i˲=ދ~DZ�t�a֠0��t��0'��h=���7�`�H\ i���FH�*�`��{M/`m乙gŻҥ+���V���U)�$a�b�p��Me�HT��/z�5IoS�L�ɶ�o86�t^xel����){�TH��Tm���+w'}��O^�Q�%��'?Dز�c�� ���tI��QşğY�v?��҇I^����h���<~��	T���U����缣���SP��wX�E��|,�̘���0:'	��K#��L���J��9t��"ܓ����.72�B๝
$������:�������r�Ǟ���Y_}F���+:�1�m	�#IrR��t�E�:(I��t�8��_ͺ-¼�˒D-�Vs��4���)�,R��2zɋ�6dO��EW�[�������:�;f����0�P��=_Q�K���e4a�P*�d`��y�oj(1�*B6����v�x���.��i^T�JZ�-!�>����_쬯���ؐ�{�h��z���Ec�v>OxKB� ڞ<��QD�?ܓ|�s hJ��Zy�m$�B��,tvx7p�ݼt~��.���?�S�\�Ŏ��8αyͅ�=v=%����R�	 ��o~�E6#\�I��ԫ���H����� ����SQ��Z}��F����:�%�=�h*��YG��S���,*� ��U;;ʂiF2靋�QOދgvyxs�=�դ��RBm�}�'Y�t��H�#X��%+PG ��1O�x6K͈�;���������Gmi7�O3�;нQu������9l��1$z�P��穭
���X!�4s
ܣ�W�|9Jk;��g�}?�e��G��Z���:�菥+H$=�4�|�
���y�{�וHJHLp m�F���N���>!�]���c>��vҮ�$;\�������q���N�s?�`�D�4Y�	���y3��U��|̘;��"JM�[LU�C
�O��dd�p��kbC�)��rQ۲�|H�vw,o���J�θ%��rb�$v|��|@x!��(�F,��6n�A�u;������Q��_?��������$B�P�y,w"�Zo^����9�[8���z�>���L�2=����T]3Ҿ.p!��Kl�)�C���Lg�\�\wTS�R���1� H����2���*�XDF���P��WJfȶ�D�F���rz�`�-i}��$q+�>%��S?(V��9c.cF��W����k�P��s(p�jH=��?������՟���ԥSM]�V�!��X~Q';E�"J�6ޥW���c���K��R�p�*�~�L
yel�*3�5���*"u�+�t��(H��*����L��?~�A5��m��ں�aR�x$P.�(���c����J����.�Lϲ�""�' �������%�[dȗd��`���v2T�$d�R�SA�d�`��w���m�雃M�uVA�E�w-�m�1F��L0Mnb@����UE�\둝�4���������[�#E��PL�4��b&�x�;G"M�L��&a�/O�J�=�ק�wD	z�C?�b*�kq=��~���]�3����9��壚�V�	 ���m�Zᖁ,\ѡ�����)���%/#�$�}'��P����a��8�eҚ�7��E�L���KY�U~z�d{T��(%7��Ӕ!�4�
��NH�nzCZ��WcX8�g<����灪�|t;>k<�D���vV��\�)7>�Sr��]>x�~"7G[�z���i^����);��%[�"�P��E�_3��e��EGn��UӼ��u�[���ݷ!��:���3k?6��݊[��M{�4Y�dY��{ſ]��띧ICM��`�PE�(���.PJK���u0.�����:+�_h�'���wq��TV^-~��s�	�SU��5�4���}�[�BY���_�)S~�۷^ jaL��	̱(u��쥜A8CbTJm��Mi���ks���e��6������k9�5	@��q '߫iV��$?4��g|��[.�4��UM�(�T�T[�=�b�;��$7���������Sܗ�����G
Z�=/���դVC���$�@N��r������X�����F�~�K4$�x��Lm�܄g��m�KS�3ga���<+��X:�d�.��>����v%�P��x��u!Yn6�5�;Xhd��>`�ɴ�~�����0A�s�^�8`�0" oQ�?������,.H9fb�s_{Ԙg�4�X�Y��;�4��.�t�h���{����ǃ%a����J���U��c��I_��O�6����*���Us{�0748�$m���E�x��$��x����{/��th�~���n��ն�_\��5W�UO7(� 5|e����^�u��+0����]����&����jn�� �`�6�r�7�}�P�{qsҨ�c��L���D6�m���{U�*���R�����TK����s�Q�`~�%��������͏�
�>����L\d��4݇�L�V��mn�O^7K��	�*�h���J���*�� :��xYN˗�����c�5�ǜ#h�U�X�����0���q�k����C���@���b���D ��Ͽ�uڼ؇��E$�~�(w�^�2q����@!6�3q�z��#HI����O�lj�� �;!��Jق��ƻ����k�������ױ^���e������[�����f<lѓB�R����y��c��AXZ�dF�ƕ�q_t��2&~�SD#����Ԃ��ڟ>���f����}��w��LF/	���{�S2-�;2sU�d�dD��~ӓK�W�aZ9;.����8wU��NO�/(����	�"���#�etgK��M�ځ�!H C�R:���Ѕ��[:�{����-_��ل#�t�����P�̸�Ô��y|w�wi�&o�~K�4��ҿښ8��>��M��Z��W��5,�&�@�a�i
R���05l�
+���6�8	�S�~2�>��.*��Ϗ��#1O�n�ۤ��vO�j��3l�t�͍����TT�~nDQ��������<��H��3#�FewU�4\�[z�.�J����4�'ˣ�D��ε������]x��,уsM��8��)9[wPh ;�S��x�i��.5eX�S�z��v=�'l��?���X�q���z�1_��]��FOT�`O0D����L.W!�ʘu��Rݺ[�s��#I���Ȼ�?,d�2ű'��A� �;�Z���`�׍~�,���|�d�b��� Y%�G�+����""�/��.E�
"�JQu�:�z0���#fф6��f~�'�ʴ'��{?��ĂX�}�U5Z�M�<�"���2�c���>��/��o�/g1����P�1���_���UCg�k8~����r�T�[G&/@�Y�rU$K����M'O�p���Wp5�3����3NoV�b�~js�T[U���&�2j��Ϭ:���U��z����1�7�1�{�/bcb�9�o�qpX�&,��1�y�Hߞ+����l��3�(��"ai[�V��3A׋钎Y�����G})a7�]���u����z1���7�L^��.�KMK���\X������sL3�{��>�=0�N��YC����3�F�w�X�܏�Gi#t������ö��F�O02p
�h�����<&���x�@è�xq=�o���e���b)Z�vs G��pLJ�$SaB�����d����a,����"�W;g��w2������x�r��ƨ�������#a�C����`���w��'��m̜���=������-���E*M���@��ի��=�t�of�o[��I3¦{�p1S��:R6U���	7�R�➉�Sd9d-S3
ƌ�@�����z���<6�shdF;����%�e3͢/.�$qwm^�~�gх-,41��ox3�gm0�jo����aİ'�f�\�^�7�}��� 3O}`2�����5���u�cׁ��:mU��x��x��;����<�.���vʒ�o���k�m�w�����>,W��G�j)#���]I������v�BS�M<�3�e}�*Ǫ��|;F�<��·ۙao�<����͇����*n��E��K�?ԗQ����#v`�s�J��	�'�����K���e'�?:&�3�kڗ�R�]�+~��%]��f|c3�5qe���3�z*s��]�Q��)ROM�4���u�A��d��e-]���R����� lR�����fhNQ�e��N��o����.��S��'f9�|:�H��,�����u�-E�(SաQ�^�_�xAL�o��8	R�.���7� %���C�i�i�B0E0bk��P�#g�S��g\`�]�+�ry\�^��V�2P%�77�lf�zZ4��eWm��e��P��+g"Z=c�
����!	wu���+��D}�|Q���Ǩ�t�؃Ƕ�<+3�Kn�Q{}���*����bP�``7�Y�"3����/n8�6C���MQT8̅;I"p�o��0�^��k��F˄�דصM-E��I���s�j��[�)&�?�o��p��,���j�fn�zV㔋�>k���fn�&�azj=���?�9�RCx�L��8�  �r[����Dg#��y���崤�K\3��q ����V�OS����j��w�;OB:���\���3ibte+��T�a����?g0�e-�y����_c}��ߩg@��©�oG��K��x@W糚>oc��z��$M�_!>�W�w����\ݸ���K|��������Ku�2r~�K��1��Wg��i���E��̅���t�X�
��`�K��ǃT�Dg����9\�;���5e޵�[�B$�_uLT���쮭���:�1Y
�y|�FF�6۸�RU�s0W/��*(��S�z��B�H�.{�SgnP�&�t��=��oE��z�8������	I�V���`gT��^@�b ��D� �J��ϙ|u%��i����7~�z��B��M�1� w�A�^V(��oN��f�A�:�����G�x�W,�D�f0�`��J�X��Z��M�(=��uO2S$�B��>X+��V������{�'�/.��O�/|�3O �=���ᜱ���)�Z�ZA�f�Ш��w���i��uu�w\nl���Na���V���&W��U�g��;��S��V�A���Vw�����r��;��G��09�:Yz��9/V̑����Q��$@#z��M���C;:�Y��C��)�m<L��)�Z�ߧMD_u-�<DРޚ�h6�0�i����h4�d��zȽ"������- ��7�?bk��i�� �>�+��ð��\��cd�Uyڮ�{�"9`V��*���X�y��޵�f|�6�e��u��	Yo�Da�YH-ݲc�;k�*e/ʞ���w��B-Ds��*V��j��LZ7h��j��>vn���d2�!����Jp�����ع�X~�iF=��M-�Oe&��gC��DZ��� Ƌ� �DV��"������x���?Kk�{

%Q�)�����@��U�����~}�EN�$���.
u�'��]�K����c]}N�ģ$����_����;U�o��>���; ���D�h�a&Q��< '��|	w���E�4s�_��f�;��I;���`�6�i[}L�q}J���z�ƹ�PlC�*?2�,Q¸G�b�U
�o�(foxp���w�O�72�^�I`�*�L�Sٓ#���A��u�D�i{W�g6U�Sv%0�R�@�����Qw�P�g� !^ĝ��l�� ��
�D@�;�Q6_)��b�����q�,��6��c��y����l2�����1˅�Q�mds��煝yh�{~*��]���e�,�_��A�p�mj��`Ҡ��	3���GmmC	�ϲ<�;J٦q)+d�wB�&�_�"��^�(���^�~��i����"�|K���p�O� ��8.�!>ny'���k_1�6������U[#�0��!K��R�� b�2Ea��L��g�5��3�I�w��o��~dI+*(�;�n���q�F؂
1.ٲ�p��p2y;p�T��@�|IO�S���/�V~�S�R�D��T����\��m̠����ag�^k�Sԫ��_�ء��^���Jm̢ϼQ̦��$P|?2�f��S����zU�2��H�<��o�Z�m�e〣a��]p�rTP
WVz6~��<��!����Yy=��@c���Ǽ,��SǸ"�䠩ι�T?^�>������}]���f����P��i�'�/j���Yz��9/�F/�@"�^�}V%�=�^9�|>�d	�w���"��J��jCM�W��t�g�l(�q�2X<u���V#E��f��E�ж��x��h�	�"���l�^�Z�sc��l�`��� �/F�<+e�!�c�=W�w6VXC�M%��g�I�A�lPkBS��쇨se"��0�؎y��N���Lk��m�/���8�
~�s�ڎ�m�	��'�`5��.��o���V|C6K=�LЪdѬу����0m@<7�T���6��b��x���o�*Ѳ�bK�)���5����Qq5Ѳ�<����nC�;!�;��Kpw���-�C����w�}��韧�쪮]��:����h��m�񹞫�z�Q}_~f��
��3z����Z�$���+P�bop�4J�؟e��[|���yv&�l����� y���Ť���GU��u4@Vت�V���kb)�OW8�t���L#������G �5Z�8{<{�%oW@����`V�n��?��@4�A9\<��h��܋v��o���^��ݹ8]��Mrl�cuV��M��{c�M����,q���J̮��!'�N%'�6x� �������pH����QtOs�2Ŝ}�$��-�Vz���R�;��������!���}�T���e���SD�-������w&O�jm�/�$T����� �T�ƛ���s�Ȇ��щ@�+~���{
R֟�f^_v;{Wm�P�9o�j����*��1t���K^͓�z1zO@�?'��Gl����Ā�&�k^�2x+ž��W
~W\޽Q�×������[5�?�|h(.�e�	�����
�;�M�r,�Akv�� ��k�iˇ cSRu�,�ߓ�s)W8�@�U�����խ_����)g�L��
'5���v/m؅�}���1�Ыw���@��YxL��i*I�Q��ڟ�U]}�n�� �B���G���;1���A/�rO��.��������_��d�!��.-I�r�����M�}����"�NrY�.�I��H}��K��[T�|�`~M��<��+�_Xkm�]��?�=q�gW�;������(���?U��=0�L�.m؆�[�����S<�a�SdE[�����}�]V�@VJ��wb��ܺ�������~�������R���ȝ3o-߆��n����,��Д��A�T4���1���~��̧q���Y����9��I��$ɖϡLߣP���p<TeHj���a�NuX]�ɷ웖��J��}�5��6$�,`הￖ$:X�#�m�������_8ڡz%D��$]�#��)�]���ng1�����������5�i���a���Q��{��P����-�ܻ�K�Bv%V#����;a�O�Q�P�7W��~;�^�) ���{.1��f�L��i��(��m�XAؘ�2�g�a�9�y+�Qof����Vl5�utG���������ބGī��(]�/�fK����m��)g���)�߈����G9���v�߷w��Ĺu-gl~����}Mz/Ϣ�Q ɓ?�p�Y�77�?�+��dj��C}����g�����'�5-a����p7��!gw�#ٖ�S�����񈚼mC�'���}��}1K2�2"	��Ns���C8�Ø�CT�ضB�J���ka�٦���W�a�K�|L�n����m�'5o9�9��8���i�e#��O<nu���Zu���̗��]�4��ɔ�`�ɖ<>�0=7bw��2�$o)o<�ɟ�{�l!��a�����a⴬[񭲅� 罦n������T=�p��^��}��G���0�_�Ox-�T�l���9M�s埿F�U��wߵR���.OB+v�}�Ѭҭ�I��$���<���E�������UU�ͯ��p� ����܆��爩[�e�8.{M
���lB%B�*���Y5��7%�	�T��ƚ�	��k��L뷛���$i��/	��L�J��L� aЎ3T6�
�k�~�D�-� SI�~1H�`"�DG�M}������7�*�T����d��׉5��j�t@D��!�����]5ș�1��M~����V�%��v�v�0*��J�,����t���'��:��7���%;l"�w�� �]�������w;�4��j|���}�N@�Y��d~��&��q�s�.�VF�N��O5*�jǗPM%V�z/�}�K��HE)��f�ʪލ�!�+���\U�K���3�
:�Z�{ձr��S4����{���%yf�y�g	t> ������4Z���pR��B٘>�~K���+�p�ޛ�6M�8$Ԙ�X�{0�q��S�8���x1$���'��5%+뢪��O5z��Q�x�H���ܟ�����һ�C��d%�r�]���/��KZ&�xqV�Y��-���m��;ҏ��?k��l���8��*K^��:5����֏syGF���Z����\�8E��.��9T��Ym8���
�B"��LnO		�v��Y64WN�B5�r8� PL�7 B��H��<�v�A�h�9��|y���h�~4���c�8�����
��Mq[����d6g��XɂeV&��2V6:6N<�p���Ԗg�l(z�Tg���[�7�M��4�D��'T��	�������aѵd�HwT����!��{qRrsSO�M���J�F����N�1�J��7����z���"�'��$aG�ʇ$�Sy줻7#���L\nd�Ȃ�����-r?�P�='�"�y"T��$��O��1��|g��w$�; }��c��J���u%M�G�8�־�6�V�O���[�<���<���e_N�Ǩ8��'�_.Es�V3`���zU�بӂ��X���f��(���g����?.u@W��yQj�)�H�H�!���������ȶ�s������tV=��3�zV�д���X�m�?�Ǚ<W��U�(Gs���il��J\[�;F�t8���]
y�y�q1��)��~�:t�$�����fXץ�0�3bx�|�e�E4�{����S�%5Is�E3� �n"�?��&�����	B�=T"��/"J���'6MF��Y�2�_Ɗ܈:J��!^�y�F��}�⤀U�3�l����u}=����"�rl�V�]j�￻T��r������ฎk�#S�����H�X_��Al,��3�5���Y���g�g����u���}*��?�g�e���<�1��)�U��3�*B�n��Q���(����=԰� �	�F0��aM�C<yS��K���ɲ�;�}����2��?>Y:�u�w��1������Vq�=>�+Vm��Hr�Ѽ������V��5���Z�<:�LR�_��K]c]�
u�͎�x?� ���/�P0i K<ѽ�IA�1��P���F�cYv]�CIǽ_(]v�O*���x[>|ؤ�t���V����rnIU������&��9�&�\:�o~�'��%VN�;#� #ȫа�)&=k��3��o��>�6��Tծ���ԡm]c����j�H��	�s�d�2���-7?���K��Q�x+��k��1�it���՛L��2CWR��p��5��G�8e�<��jϑs<�ӕYS��*�����7/�ǭ�<)�'���{�Ur	�ݣ�v��_;��� ��M�q.s�ߴ�]8���@,�^�ZL����9ɒ�h]c-ac��>iCw�bs��W�ņ�* Zo�l�{A�FրN7L��`�~[ֱ_t�}��?�6pR*]ӳS�9Yq	�ӂg��G����C���et�@�
�����I���!��{�_�U��V��dN��\*}F�Z����FȜ�:s��H�G�d�e��>�EWN=�=��n�c���)��b���$7wxrC�~�Fz
�J���C~Ϩ�g��@k}8�f��^ /Qy��<��pIiK6��I�[4�
�5��m�>�Y���N���l���'U�Џ.��u)�H��F�>�2��y2�[�qjn&�հ�\���b0���~q ��1���
A�����m}>O����-6�6�����i�]+�~��哞��2x�� �-�Q.}�KW�.0���ϫG�Ivu��j� �n��0TP,�<�5~ǳW�HW׎H���K��%�sS�e�z�0�LP��0��ۃ��9񛒀�#�Za��<2����05�iˠ>I�m��\�7�k�&��#1��u�.�� "�~�/�b|���ݟ�� *���1r��Lͪ:��E��$'/<�,��s2\�����7*� 4#��hO	�r?�B�Ή� �P]1f@���-�p�����]9>UL�,_7��"Z�E���.�n{k�P�fi���ۙ���\���(D 4�M�4X6�'����Lz�Zeƈˆ#��[!����������@I�d\����؇`��e�>�aJm������0vՏqj���ͽG����.�&O��`�'��'�aY3�����P `aV��n���pV��O<�v[	�AA�R}f�����G��zN���
�I�r�[	)h[%Ihp��	V����+COW��[n��NL�E|��Xo���0��ԗ��i��HǙ��a�=��w�E�Puп��}�^-�>�%�N��O�>��Z[ Q��BJ��A��]4v�+ȝ��S�k����j���dJ_a���	���p����Z_�%���ꤔ�#���HM��s�'a�C������W۝�ot�ߦb �	�Z���tk^�ܴ�c��	V*V�?oS�������58�I�P�I& P��M�q� f��R��/�z�ͧ+�#=Q���@�����
�k��a:����������������r�dBɭ��TD���VՒO5����s1�����{�ȒB�j���ț���a�:�7�&��/����S#�>ɢ����-�	6��g��I3\�%�x��"�5����S�2�x?�lMAD�N8�Eh��8�Q���r~��>U��>��Jˇ����;���YF7�����
�@Ll&���%2���[1�V�f��!�}����9����(W����c�V%�����h�����6�夙A)���
?q&бeuy��?u*Ԗ��T��Ե��b��"W�g(!�9]�_9]�V�64���E����f��a~�������"}�q4"����H�d�d�MYlT��B�}�F��(I�`�F�2a���tP�c�2.\/z����pL93K�v`M[����DJ9cL����)SQW�@�^�-�1}��	�sC�$ �\<�IO�#�+�$]o�Y,��ۡ)Z̷�
T�#�d�˶��";�����_x;{DMU̗̍�Q5���7�ZYȚ#q�l!Ui�������=�ѝ��YE��
�:���@�������f�G�n��^$�<��g��p�k��Xj"�W�N45�� `^j�}m�]���\]��Qt�^������G��f�x����� ����.�*��I�^u�,�� ����F�R�=�'����w�h���'1�z�{��i����q�DxA�`��@L��.O�6s&�m=���Q�����H������kQ����H)krM��	���}@��3@{�^��J9�Z�3�F�=��>0�Б�D7YJ^_̼z���?4E4�������^�w|A�^=&Du�R��s[K���D���v��.r}�� ��-�U��1��qz��������{��Jx���Q&�i4~�8��dr1b�H��fS%Ai�En~Z�i�F���cE�m��[_�W+��BQ�5R��v��O�{��n7���P�y�3�rɷ��U���9K�(�R����+��l��T9p�_u�g�ʅ�q b������d� 4���]r͂r��H���m	)�i5�qe�Τ�Y�{%�u�#4o�T��3� O+>P��-�x���9��Į2�s�~BӼ(Zu����-�K�f����s=��f�ӡ*�������IV���&*���g���K�V�QR(�r������ix]C�q���Q���h��I.�eL�*G����4��k�+���I�p=�}����mW��T���?IT��/`%c��o�,����5���n����(Z����{9��٫o����E�R�nL"��d�>�:��e��&{T�jh���Y-F4���t�"�s�����	�������K�P���Sf��g��I�����ھ:)�Oev�=��,������ΰ���.���Uط$ fU��R�zVI���W�-u���aZg��Jb����6��\TN��%E�0M=Ӄ�q^H�)+8פ���D���>E���ؾ�l�}��z鹬>a�Ml}�1�w��S�#>��o)�����,��3�@ŕ��(�C�!�!_�ЈT�r�Y��W�W���0�hfT`6#��$SGm��KM�5��&�a���×�����T����;
��ԕ ^��rY����*��׵���xM-��j#��w�c�쫤{0Bq���i���̱�)�a3�A��m=�r<P�k�o��g���,찭d�렽tc{0��5UO�̪���q
���$�.-!�<М ,{Qr0�Z���6�]ϜK^���brA8<V�B��3/C����t9��v�W�����V�ׁJ`b�&�Be�UY�0�����/���;^�]Pv���{�ɦ�D��i���������eh�x$��T�k�����T|�Ez픃`��tn�%��}��Ef9�hW�F�)˯~5�`��o�r�K��|.i~訕QՈ�� !�#�H�c�YZ3������]���� �F�����[[y=b!3�^��f���C�^���#���{�����_��9l9�s%L�G�y?J��̜�:�rw1_��R�·�i2.����N��btI��WX$j�) ��փ�+W��A��3��j�A�a���,��%�<(��,	KMV�'���#G{�7Fj�p�`q�����ng5A�"���ש���L���ZV��^ePe���4Զ�O�E&5�i������}��.Nb;d�����eP���i&0͚���W�<~��Y �y��Ur|~z�ۯ�0���9q+`�[��nb��>FSS�ł����B]w��/�w�����K���yL���m���$�bI6v�Q�J���x�g�t3����Y��� �QZV��K���]B��~�������r^1�w���sx�v���|4&�S����Ϧ�~�c�+LH%��Ւ����Bo��uy�����i��8e�R�F�hĐd����G�.��^��)�lgڞ��<o�a�>�^i{u�������#���(uŵp��f�˲n3��N����\��Xw������ia8m����W� 痜��o2�V���յ[ Gfm�EZ��g���(��p�NosFDd de ����A��h4�"ӏޟPE��F����~&T�7!A'U��6�a�v�*OZ�Pvĳ�:�u�l�N���I(����13�3k�p}�=��U��u��B9N�����jG���㍸or��"��Н�Q��� (7=r�9�(�-�K!�ٓ���ZO���vx|B�ψf�_��<������AA8��X�ęU���y�;ت0�s���ma���O��M�%�� @rR%���l�6>��M1*�_"�4Tx���b xE�Ek?w^�;�;�kz�,�Mly����4+0�l<,��(B�l�9�?|7E�F�+2�9�sX4k�(.�ᤓ]U,h��pխ�A�� �7���څ�N�l��kE:�Х�G K�δ��e�db�߿����+m�׳�P��ҕp͒��6�EG�����G���K��D���a{��_�6���j䴵A 8[�J���m�}�Os��O.�wf�������^�٥�+��k �hO����3��S��飸W
%��s��> �k���gTp嗴t\SN[��܆����R�o��F�R��$�T�~v���>S�?5?��b����.��a��������u6���G�
�Y]	ELh�]�I�ﻊ�7ĽD3�>�}ivX��
b�����U� �9ס��p��06�whC�l��v0�W��F��{Zs�7�G�]F��'��eY���;�kp�"����v�T=P���hg�=X>�(m�#�w�D�yi���/e��:�5�z����^ç�\� ���f V���t=}�Tb��<~�����o ���M�Y�� �, �z���h����0�.^��D6FIA�,�x؋�8�*��%X5��1ݵ�K �.f
0{@����P�@�g��-��N�|Ƹ�:v���9�3X��k��d�bQ�P����r��8:�$�rQLH���|�`]���Ud� Al�X^�ں]�x�~��>���+B���q� NyTZD\+n/_��ry�� ��/`���i�?yS݌�-Yu�:v�g�aS��,:)w��*P�`/��ho�H"�':t[/a�W�z�����;��lk�cFO��୛RAH!��.e�?�7h�[V
Xg�K(kB�:}~��hv���W��B�t�c����˘�ˠ���g^���G�6OJB�|t�u�_L�G� ��WS\�
�|���˲M�<�Y���( ّ{b�����fq�f>
,�	O6k��X������ɥ�Ni��� �E6
,���:OA
���q�x�c+A�0U��8����V�ʉ"�����d�ns�U!�Fa��Ou�D����q���仈]� �h�o�|��`�gg@J,�eo�l�T53���oE������f.�Z<�Yݠ�F~�U�#�z��sثlN��� +D
	t]��a���.PO/��)P7MR����A@�Th��G��xX��'>E��v� ��3�.Q
�/��i�4$&�l��Q��"�J��kS�,�w��U\8s�;�C��v�0����>�X~� q�n�:_�3H	��L��U.�,B��:4,�j�!�2(/�xd�`�I�[����E�t=]����H�`/�7��'���n}k�����7|����گo_�J�Rd����?7�रЗF�YP�7@+�_�^�g��]�74;Ep�+�p+���xH�����%�Ңv9��������=ޜ� j����k�A���39���c�u����q��94��X��H+��Ъ�OV���ng���������#�7T�L�*t]0�P�X�\����h��8��ǡ��E���^��m�{���2߭��AD��(Ȅ#�U���au#����ϭ���)t���:���e:�IZ<�Oh
��Q�:j�u$��ɾ��F�a�ظ!!Cd-E;�Byh����1��c���o���4r��R�� bv��C������A�^�RE� c|�q����;}@��t.�mWć�6T4��)�,|!��ٙr�|�� ~)0t�_��Y.�G
 ���"����sOxc�o�+��&�rTN��^���ِ-H@�Ja&z����3*�`�nd�*}��	n[��!��XeE��Шl-�m�5��T�.d�={߂�t���R��F�`_a���&za3��������8*A��4��.�_���Q�H�o @�]e�@�Y?��%�U�%��+��Ƚ�E.E8���;y�����>4,ܮ�_��(.$ v�\$Ż���I��h"�CÈ,�  ݤ7�Q7�ztI:@^����`�&��Ž}��/��Q���a��*��b�G�!-�H��Ʌ���03@�(��Q��������6�߀b�oF��D^^7�ż&�hDD�E��D���	.k����5�	#�h���n�1w��Om�NzT�?�t��R�a��#�F��n'=qM�!��gmk�#�\�ԒPpr�$�U�>9���*O,�*�������IǕ�Ҫl��%�.���ņw��(
z�c���iZ�Qu�[�^:�<�ዹO��.di��O��'v�`����Z]�a�Kv
 h�0)����^��AB���Ә��9��=cX,ꢱ� �Z����Xss�����a��_	k5���  ���!c���y?�F������[)򸟧�H���?�����+����	؁I�xi���rH**Q�A�'��# 	�+8����w�G=�Ucoofa��������	6g𵗾	;����g�7�Ϟ��IӘ\�ʝO�{j�
b�Q�*9���-�k�~��I��|��|?˞�Z���>!ؤ,iEf��ތ4<�,T���a��\M�J2�K����jٺC�V%ŜI���U����F�c�#�Z��P��~�^�P�R�≔=݇��Ǉ���ɐ;(�k�^�t���v�����_%�d/�
�J���>ܤdH��#K����ϓ5EǛ���|��wL�e�^�.�k-�Z���d�?
���E�i5L��.��M�lgw�c?�sS릂Ɏs��2��+��U���ʛ���x�P;^2N�B�ܔ�D�����ޯ픿n�������x귴R�� ?��u6��۞�;~y�����Xq�d�W{?��:���x���^벆5���0UK�g3)��J�{G2@1�ݣ�"�Me�_s���4�����u8,�]���F֌��=�}�0W�
�鹳 2�������zX%�徸�z���h��i%[��%t�)��� )�k˴X׹�|���.�n���c���=�u�����@�m��Կ����֭(��[V*=��kU0��_'���/������T��"���Bt�<���y�M�u�2,�x��X
ƽf�>��~��3Ӊ�m�X�Uuutސ�����>=]�I�L�� �B���8d�W,�2�k�G,H}c"j�I9pdO 0���D�����>e�4�M%����$�~,��,�k%:vc1��=�����Ĳ�̶�y�!$�������ۆ?��F;��H1DL����d +I<���s��t�l�b���
֚B� �φ�.�	Z�O����}�2h�vE�M�<�Zn���M�zॖ���>�?T���kI#Q�0�i�okIs�{�Sʛ}1N��W o��7�ff�ث�}���?��U�k���=�d��[� ��rJ(�E���|�!��Y0m#���e)D�Κ#�G�Ɖ���g�XM�b�&X�dÆ�]� ���!U7x��b�,��������\�� R�]�܋>�`w�c&'c ��_�y�M��ɥ�Ŵ�����m�J/WR# MW�����~������>��#���(�����I��Aз�=y�0mYGb㽉��"8W�
A5EsUH�j����P����dH���N���u�b��}E.[�^@��O��\��{���vVtԤ�p �}��2pO�YK�yF���g�}1fj@UtbcF����������Ռ����C؎�>"0��3�d�
��Ӆ���#U+@��3V
 �旦�^�{�y���� �
v�B��w P 8�h@b � uE mO$9]�n䷿�T�zf��sѾ�;
�aǂ�3�N��\)���<z�N� ��1a�A�A ̧̂)?0��������e���U�A-���m��`C�-C���b��,�9z��Ұ��R�'xL��:��.�_�I68u���`V#g��ʛq���L �Iz����+2$���`&Ѝ�0����[s#���l��%�#�+ kZP�"Je�'����d�m݇	j�B�<FӓBG���~)�Ѿgɟ�I9�8m�M�B�������ɢAH�h�H�n2S@!n��<�$�j&Cy ,@����#@�?����0^|�0%5�*�Oj���i+����a� �J��vȻ�5N|�"b�s�	�q��g�4tT|� ��/�4iɨ�-v0�Q�������8�Q�<�(�GTn�����{���V)MJD�~ ��]�����d���]68R��)i�_�7`Ȉ*
�ڍ� QB��]�
�Ĥ�ʣ�j��J_C7��`�Q糖"��A�!�j	���F䥀�r�JR�T׷2b� cv��"����q{�`��wJ�^�y���UQ��hK��v;eX�G���;nlD�0`:��BpO��	��|y�GTg��[�"�m�wӻ�t}�v�G�ԓ�v��_.��Y�	_��YB�0W�(t w�d�t�DO�-�ʖ1[���j'��;� 3��D�l��l��y#���&�H�C�N2��{7Y�a�)@)ȶ�!R}X�o�������O|:��=�v#��uV�Ss{B�Q�H����տ������
__Ϗ��
�8o���j�`--��� ⫓|=]����S�z)�ЫO����Q9$ӂ����)��s�"͎ �A�����G=2ߟ#�١��T���-n�l����=}x*�X�8b�bY�0�im�i�O�
�Ȭ�{�@�0{@�a��28?P��]}`�3�c�� ��5�>EBSӽ4xQ]졽;��g�}^J��;0��҈����6�2�)��]$���@R�IGe���w��%g�&��:'b�)R���T
�3�3u,�sn+k'VZ�㞼��mhv�����j萘o�b&�~�fdF!-nR�'��`����s÷�;��YJ9wp��ݦ￫�������
%�Z�W�H([׸�\x��{�k��<-4�l�ӵ��_��8׻�o)�BO!_��@��kU��tD́�Sa�xD 	Q&ɍ@��������7���0��Ί����|���B6���Q>�yd��;��.zs|���P�-@j�!�/V���9���$Z}`x,Ӕ.�t�	5�������I�$���k����2�m�9�Q��o����h'QH���0�5�6E�S�"H6vp�a��-X5`BHF��n����ᱎeiL���｟�D9�e)hM���|N�L4���>es�Xgog����"!�j�H(]\>)��r���,�8�.#]4�L3���������?�,��5����vTWXL1��H�[�.#�@�?u��6M�ۮ���@E���}�s!<#hP7a6b����5�*�����C9�N�th��"�$_=د+�u��k�l�n��ʾ�8�2\���ǧ��$���o�%D`�xw�v�@eh���t����7ؾKE�U感�.w�&��w�uyJ��S�X;��~H�ʢ��&�>�Q� ad�p.j��^��;�~�\�빾�뤔�m�RO�G�.����*��F<�	��ٺ�,�,6�h����8��1�bu�Q�������-q͉X�C�M�ƣ�B���:;GG!�CNV$�4A5������*�p`?A����^����9ן��ͼ�+��@6���qX��4��栰����@(��W%2�PhJ9r-(��V�k<�q$��,V�Όu5���� :�Z����5��r�)1M\_	�t� ���u}��閆����9҃
O��\�ux�T�q��zRQ���Kh=+�\х��%@0����;v|oQbX(��i[��f\?�������C�h���Ğ�f��w�����Z�w�	��Ԟ	Q �
V��2_>���_���
���K-)�Ko�*�����JM�$2���Az��;��Uvs(��ڴA���5��%��r�@r(xzg��D[�QG'3�{@�2h	�A�<�J!����6�.匹���o�����${ox]VZ��kM��6�s��3a����UG#�_�m�DÞ���{��� �����Ǉ�@,���<�w�1¶ޓ*� 	Iy��w���Ul#�@{p�������&���e�o�]\����VK��<dXX
x���K��(��C��;?4�&v����#|0�v������,�O�k*��h��p�L��"�_�kb#f���K(�~�j!`�[w��F�\f�o[.y G��鏹�W�l|�'
}��O�G��9�Щv�Rb9��n�7�U~,0�̆�&���nF�J��u����u�<��|��K��Zm��vxJ��3����p Y�H���)1ޕ���B������
j�g�]�j��\Wχ3"S���C��"��,	�'G����Рkj�������q���Zo�&�w\"��CS�W�(���=��Ä	�aJ�FB���X�Pv� gb���1� .��#�VK$��~xx�&�
�����<%��aH�Y
�qӂt�1XZ���/sɨ9���߭��N&`��`�^���$�\� ʑ��"�c�(���Q��݃\�Ǣ��7���:��fi�CN۞ؽAl=P���e}?5�l	f:z�N�u�DO���MYVVB`�hg����_�W��U?%@���>'0u!�٫�k��i��������#hW5։z8���0��!�&�pV'��B����(�����ft>���{��C�,wQ7�aE���]��j2υ�΍?���V��C_��ز���Ƚ�_�����^�`~֌������Y6Z�A�|�m`�{a���t�9�m^�]։�3J��" �h�����(�9���#I`Ywb��D��_2��{y~�#�سQ��ί�R�BV���E�ث�̴�͊7zMe#S\�4�H����/p�+b���� �1�b���A*�Av��Fy�G���یe���XF�ߐ�T�Mvѻă�s,�@���S�W{a+��|���X��Y��A�.���u(�c�q�xJØO��D"BTF2�H�3��19#g6�����}�ӵ߶�!v�W�]f>�:ټXj:��ۥ��� +�l�k݃�# H�9���p�坾��p5v����fM��?�ڰFv�^��G�{N�,��e-�
�]�hO�y��adq��a�_=��Q@���%�+{�m��~���|n��r�4E��P�;պssݚ��	ɞ�br�u��#����og�a��C���̟�憒�iO?v�&��u>��e��ֵ L�ﴹ��ҥ����6c.2��$�G麃�S����Ǚ��C]g�o�l��n"{)��a�FE  |wXk�)1�o�����#��p��b��U�*�B{ԗ�>�q��N��W��7�5:[w����M�e5� �R�׷�U���ܾ�K�f"V��b� �C@�j�R��?�J�?���Ȭ=�/�v�=��o���
��?t
���F�}vD�IoAlqi��Ѥun��3<۷�Ȝ�#蟭T�����VZ�
0�@���� ��%�}Lt(ِC��4��T�Z.�{R_&_��-c����O��m�򤌼��}|�_�9پ-q��ׂ9�|M ��j�,`����ᆸ���2�9gn�EK���g��՘]o3|c$D!��M�%�L��<KC�J�Z�
�/<���aT��l�n���[2�2�m�QJ��V�d8�p���%�yXK��W�/����Fs@��P9�Ma�}%Oxc�����.�U%�;V�\:m�4�u�;sO/=fvG��[��Z��T(M6' �  &e��ӊCԝ}������{���V�o-��aOA���ԓ�8P�r�1:��?�d?�M�� ���qHfY��D�����j��6�C#�韍�[�#�A󄓓z���]n- O�U�Y�sE�@>0%.��|�5f�0�t���k���m*ߦ��#<+1�d�}J�;�Q�53�X��k|���M]������x7~��5�3C��X��<��7�~�0�& )�I�#�������)��@nF�|;�r�w�ķ�"X��W��7ԯ#n��*�CSWt �K�a�r�}$�5�(�oʂ�&�&z�i&xr�h����\r�GgD-��Ǥ�uV����#�����@�W:��O��x�U��jMN�t�?��f�s�o�4��aꂧ
�	v�Wވ='���>�Jp��V��j�ը��eT�!�$Yba�T>-�]e&���Qyݒ�I<;*��J�(��m��&�<�E<Hs��_��{0�i'y�nuc�|����q�p�U���\�oZo(00��%	{�DW��fV:ao��ZY��S\3�ئ��j v�u��pG=VT��L�\����SJ(�.��e�j�3G��t�������
=����_�C���\4zem�'Ae����@d�Z���n�#,`;|H
N�u&�\��BTt�K��q�t�'��W5��V����6�a%o`u]��#iԚ���\��?�>t�y�	��#:y~al�iAUj�j��v�C����c�iR,Vg��T�r�� 3H�|���낺�(��[0�!���^D�����9�3ʗj��P$?ũ�Y!�R&�$r#>��OQG��fYA �MR!@Bb��\\�`�?{FHm8p"�z�n�/�5HE	5x7�g�꼽�$��A�W�q�N���MVƖ�b�"�I�G��)&i���o����#ri�����{�����!�o���~����W]PR���N��o�R�ve7��m`�D$�7��mϔ�e������J����~h��@���t�2As)j�ڬ�WsQ{��}}��p��Cz!�����P�a,��w�Mt�^�R��3��>���P`����E��D^�-D���]��J���~�o��Pc�Ry%ʶ��c=>����Z�,��sT>ff��L �p�3�L�\-���o0��U��@gJ��J�q��x8��:ڨ���֎��;�m�j�&il[;���h�6[Mc'��9���k����{�=k���z��nQ����?�[_�J����S4oQ.��t�q����з$s��y�=��8˓̀Ͳ��QĢ�w���
�X��M]R�N�}&X�"��[�I��՛}�[
��?�P�T�*���>p����<�,� �$+��4+�"���7`��Ǫ��<8��&A�Kꢙ3����Jd�h��Rn��i�eI������oϹM�"4Նu��6ND�0v�f`�٪J��;�7)A�O��Tb�涉v_��������k{ՙv5J=5��C��˴3���#��Ǒ�5�!�7=?_�b�\4�аٛ�qs�y�د dMO���A*sJ�[l	˘�Cŵ�i�T����!�[��R�}�#-�q�{�L9"7�_�H���L�8�H�4'T���)��_���2D��4
���o��7�L꿵D}��D'M?�*������I�5�*�Y��%�����fS�dt���xqy�،��mτ~���*���ʹH����Z�1�nq~��I��W	�tr�ے���f�*�>P�/3�SA�e��O�j�k'qj�s����h���^7� ��4�6�2��.%�S���fPj4V��IŬ)gJ�{+�4+ۡ#Q'�[5K�@{eP*<T|j�7F�u���b,�e�)I7-A��Au�fc�����I���>ie�l�������׫���u�KU����w���B'_��m
�r���f�tZ�djQ��5�D�C�����O7�:?�O�ZH�K����Wδ�q�#h�i�[����B�*�ӫ��n���&-H4��=���M��������r�;��{�d�mćM �����da�p�);mSuSal���R��{��@�x����o�\�'������>��|����,�#W6gn�rѥ�&p�& �1����<�g;��J38�G��Lm�Y*{N4+BB`)@�OI$K��X�[^�����!����6�V�����6lS��ttkC��� {�.�$�J�O��\��d�����h��V ���F� �4��c��^��I����G�eL���&ON�a�*Y�Ca^1���=��x��!S4�c�y��c���VG˫���Tc6����gJ}��6�wt����X��Z��_b���^5ۍ��S��K|��*�[E���=p{e<g�r}�G����g�@����۞j�w��T�*�@�Z���_��
'��gk[HKC#��SE[SEGS P0�9?4�=jﮆ��a%٘$��(�{�d4'gtGC������:C������?�X�;=`�ĥ^ń�j�9�Q���:7s�R)�����ߢ�b�z��\�)��b	FPQ)��Qri��b���~��rU�-�8��}�y�e�}r�Y�x�.x�+�;	��׵���wjm:~qO �c�̈N1L>�'t�+r3E��QZ�Y�"�~��U2�A77?�ځ��8�˿ZA�[��t�#�"�q��G
 %҃a��a�bp��k��9�P�_�W��2���Y]���QGc�&���(	��s�n>�(��Cj�Փ��ΥD|ȕ�Z+Y"9�U��c\I�Lf-򤕎Yg�o&;)S�Q\�Z����}6���D�9��Qu!���JQ�����"�ȋŅz�W���<�K��ND������V��W�B�	������/�������F�O�=���<h�d�������Dw]�p&��l���J:��5�IşdL&���)�:M��3!?��hU��[8(�ۏk��?
�;�:��`�tƩ�س�8�uVӇX㽛��7m�	�lm��BF#B�'F���ǵd�Iu�z���:��iX�8�Jl�Y��iw|�눘*�w��G٤E�5~�q`��d$�}�dSNTh�O�3>�l&fX�-Z,c!s*ĉ�3"$3o.����k;G�:�'�F����)�.?�����K�o�'�I�S(Wr�,����DlT=V��U�,D�w�W�d��jL���7D4%�
�V�J���G�1�N綄��x��w��"���q���f��t�d��tj�_|>�Yh�Z��>Ck��B:?[�r�� �ܡզRC9�\*zZ}	�d"C��F�,�"�B���qf��C�T�>��Qu'�6
GP��^�y��/���.�i��=���9���w>b�,j |pa���j��� ���U��4�.��2p��k]Ħ[vI�o\��B����SQ���-ø+V���+IK���k�q��q�=����剮�oS�[����|�1}\愘z��)#Jj��Y&����6K%��@qH`�3��j[�>��5J�Tmy��WE��Ļ9�������+lW�{CD�(��T�Z4l偧T)6Z�ԫ�qgGچ(<1�<�
�R�u�x����]֛[+Oڹ�e��ui&vo�]�NsO��"rN���k�� � ¿q�i؏� �k|��5��6��+w`�L?��'^���-�IGa⛬R+4��
�9�D�\�{CHI��S7����`U�ޒ�}��RS� �f
=c�M��֛${a�J� N��6<��DvQ>�Q��ՋRe@���I�2�m���o�%��1Pa�hG�gN2���>ih�q��=�Y��3��[)�&�I1���ς��X�,�A�"����yۡ�î�Ɩz~kʛ��1���7ij�L\g�!�I��NDxk�h�Zse�
՝�-҅P�S��&WP���b���g@s���B�<}z�;Y�c+�1�}f~���L��J�^+�XJuX6�^F�.g�rg~�����x�.<i>��A���M�q7���=[:U�UV�j��7+�@I����Ow*g�w9�9�HNV��9|U��E����y�:Bw� lխaҐ�6kk<@��Wۼj���t|��ex��+��DD��S'����#|=�/�䐶�hg�g(��T��W�ʴq�J �n��h���>��x�{(���F����p�p<c�M��p�7!t��d��R�h?(���\��s�cC��lr4@v��K��X`Lr���ĵ����JǄ�����>�F�h�wc@����-��&���3n:�[��'&/&��v��s��Q��[)�F���+�8�[�kqAu�
�*�a�#~�7D���3e���T�`��<��^���*H�F����R�N�m�;���WX���0"i0����6r����"�jE�{V�� ��r�.���:BQ�K�������j3��w�+�Vw��ʉ^FK�.E������;����S�t ,�SXl��徹��
-E]�7���A����Wr\�ѬNJo�C��3t2�ymh��\}�W�X&�^���q�4vC5=��O:�p�v�u�3�R�\��P#<%�U.�]H�rT��:;+�hH``����	�&�{��Q �L��$�Ǝ
v۬��a�L�3�c����'�,��;�犪M���h$�`�|r���B�	\����>ʀWc]�TKtm�<v�� �^&�ΖZ:�N���yiʊ���D�r�p���HUYdH��,"1��N/�$�D ��`ʟ�D�&�x��&�i�7)�@
z݀ϭ��
;�e,D��34�v*���8t�.�%���(�xv�R�4D�h�%B��mN?c���#;p6���G���]���c�4!��m'.�#(O���"�<i���-�f�������c��e�W���֮�ǻ��^w|��߈{���SU�-���>���R��].x����[�&�a\-"��'cV�С�+<�H(�Z�����Ǝ�ϑ���;�{S����q���oM%=l�/�r/���nﰖHT�M=x���`�vô��?�B�����<W<�[���*It�l']�Rpae�ƥ3R��̛��^�������K��#҄WO�����[(YТw����]rU��3����;]x
W6�	};�w���ٻt���5��¶��*E
�sd)>-���6脕Z1�zKI8�RD�K,���h���{�*��C��ޙ�s�"V�u�
	���5��z�v����ײ�f<g3a�B�������Jsp�T��x��T=�ݤyj<sm91��7��7��x˷�CD�#�JW(�XA��zo�I%�a�ߡ�4�u�R�?�����Ĥ�ͳa�Λ_���R�/1t|���`�4,,�e�,���a
/�5�����=m���V�%$���	���d�ɧ���(P����ʐ����w����rU���q��¦�-��Q�kp�]�򟢹;$V��r!vM�貁���mYIv�&5��A����'͐�p���0T"lVu�$���ɸf+H�.6�sv�d)P���5��>{xm�^1ED��a�V��ۢ�-ٖ�^�a���:M�č�����&��tr�ő5���:���i�D^aU�2��;M3�hy�i��3��E2O1��}��RP��g������gʘU�iy�
B�� ��aĚ��p,ȋ/�ݛsO������y��ի"�����\���-Χj��g')T�X#���,"�w�?��gZ�����P��<юh����J�G�?v`0h�+\k�!�u�~gS��8:��B��/Qr��-����3����7����Kum�Iv=��H�o�ܴ�l���cJ�PR�W��Fo��)v�;' ���1ь�܌���#��/����hS�b�,'�p�E�u��6������	i g�xF�p��F���,>�!:H� ?+�C(R�)�g	�vȥ�za����Bϓ��UG/eڗb.ļz�i�Bc׸�h�0q̛A=/�C��6'V����|CK&�X���;|; D�C����萨ys�hk�W�&���R����|�,�F�e0�<M�~{!M�EYT�`��2K`"�w(g<�:k*�7�c�@���6}g�\������Y��I�I�^q�R���
�grC0k00��_�QMk�Ul�z���J��i@A.R���"��t��~��s�*���N.L��띰	l��@	d��
lly�T�{V�pBY�z&���
C�+͎��T��cE�~��>���R�1��PY�T�~�$#�o��B��>ߜj} �&>ȳ4	�=��If��[�Uۤ=b���P@.��5�K�	�-_❙�cm���j�'tdm1���rJ�3 V�����x���I��UW0�!ñ��؊����FH���������媥�>�s�q����܂��~n��_Hu%	,ɚ�
d%�y�-ȧ����:~ۻ������ �Y�@�rñ�[��{n�"(��qP�%$��Z#�����4F�53��w�k_2��j�^W΄`t�dPQ��oS ��KyRέ8��kI�ns1E��4�>C(M�������_����G/@]��P�k~}�گ���N��T��q����u�rKۮ�� ya�C�bS��8��������}ѳL��e�����Z}s��.�e>�ϗg��P���K�--4����e�5�y�"Us����[�(H8e��Y����+�~�< 2'�������U�q���';_쨃�P�#ⶠq���A�(��x�m���V�����b�x����o6��Cw�D֌��~�"���^{���LcҠ���c�`V&[^�#������y���h�M��S�c��գ��
m�R$�}�ǝbW�	���}��<�iH�'�|��-M�vq�Q|n��p�fK��ކ�|7��0<' h�#he��7'��r%T<��.N@qj��*[�G ehب�U���mH��0��!����
3�����y!����$�mV���]��.���G�4+d��5�AD&���?+�Ts�1ʂ���V�M bi6�����y�;a�z�S��qW����u#�I�kt����Zxv��j���ۛ��B�/KH	�?���3~�P{}�+���vu��)v�v�iZ*��[��*��y�^�g)��3�,��}�Y�E
�p�uvUC�d2��~�z�ʓ�=� �Qa_7�S6���t���$�%���0�.���yᯙ�Ƒ�"E&�pPA�ȖW"�?[΍��j��0��f|(+ʼ[��m\Uܼ�(��uS�UXЌ
:rD�"D^3n#E�9��ٗ�x<>�VD�{x7=�Z��p��X��ۋ��l)T̈́�?�wuA��������i�f�Ɉ�����q �'o���@e�(��J)Q��M�숾;�*�5'~�I�����:��)ut��re� NCݦ���.-4$��B����� �=�>�N������RYӔh��f�]-
>��nh\����c�/��6\@B[SKN -��q*g��[lj�$T͂30lF��d�+I�?6�-|A�8��T�\�A�\�n�p��q�28��~Ms�
BK���o��('���ɗ�H���������)2n'~�]��.4�(	2�)�ʦ���n�:�����k��H��=�e����~�2����{����?�mV��3�����N��G���\�KL��X*^���e����}���7�Ⱥ�Oh���T%��� �mN�n�p�z�S�� �*�<�¿UǈK޻Ϧ�vڦ��̧C��jU9n,���T�n�H�����9�+�.+�>ט݄�|L뻓܌��ʥ��>���$�lP�T8��a��:�����D^�>ϐ���}�Ry�2 <ZOť8L�$��P
�$l�b��`�L�u8R�Zk�}i^<����^4N՗j�1��}�@9��j��W]��|:3�����]ߧ#�M� �I�S�7,��{�}2��<��W�wcW��T�"��.�O��U)�4I���?u�t��^�Y�&N�)�cY�EM���ƍ��(l�!��
�6!ʵ=8�*��
���]Ԑ"5J:�@RbC:���z>�Ž�;��\,ń� ��EV��u�O���ZJ6���r�%��_�I
�����+ƐJ�����6Nulao�޹������G�>��ة�!\U%�t�����n�! hLZ����4@|wU����n.�i-\�xE���&�R�I�����ѝ���Q������U,�VC���fW�?]�^������x:��_�����|Ɣ�5�>>�x�8�ւs�31V�D&'�����op���r(����c����1فҒ�+s���HlR�G|�y���bKhP�;?΀�^�s��$�<k�݁�����������S�Ʉ�[��&p5��b��a�߁j眞%��Cp�K�$G��`ΐ��.�4,2$�e����FDJ��x;�Kqw|%�Q��Soc�Pr��.��q|�y9���|{�6��'�# �vI��E:�d�;�`r�y�s����㙔��-o�hYB9�OQ�/��&���d���@Rd�:4�n8&�|	@�]���ȤY.�7�m��"\&��˰�sk6�����:�>�&��	-�A��"�_Rʎ�d���Y=q
ax�� �����C�2b�`i�/���l��P��Fv��`Q����D ��65��,sF.�t^�����='������gg�J��d9l�Y)���u����v��y�	�ۙ�@����Qb"W�h�A���v��=��$�	\�N���Sd��ף�e�V�/#B����x7�g����Gen�.n��Y3��E�1���]�`�T&�Ͻ�6���R��p�.I� �1g���h�
�T��Ϗwǫ-?(5~"����7v�7`��e�8voBtO���
�U�ϫ��W�����cۢ�C�	���!�nmɋky>\|���"���t=��Sf$l���@!���EKt�Pu���'�C�=�E0)i�0;�g�ł��D��bN�1�M����j�Ͱ��˹�d�
���OSP&¢d�>�H��|��P��-��P�4��8�Z�����n'[}ˮt��K���bBC@�{\�����
�ߩ�v�n�3������)��d53)�(��F�G�M��`#���{�2I��\>	&(ؼ\B� �|~l-�DGD4��82#����R�ğ�j�GH� 愉c�c���9�;0f�7�#��K����.Tsd�Əh4dYV�>���.��[O��
�Rz(�-��'��?�Rtɡ��W��bҟ�V��9�@	��MгW��e�T*�D ������g��c�;���M��$` 2)���r,�!Z 8~@�Q�K6<][��x�\.�8��\__�������+>%^A�)�m��?~C-5⦉l�0Wҙ�7� �Y3����z���� ˕�&Lmj���bL���ewnȥ�6�^݃��q�R��aT�oE��#�+����U�8w����ܷڏj�D9SH
n���H -T���I2�A��SjPG�پ�������~|��>�_��X�H�4}�;��F4��w{:)��/!�Z5��sru�����(+!�����@5��$+��~�=.�����@5�D����j�����}��D䇐�d(�C��'E��V�:c�l}G_a��:�x�R(0���c�
��Y�0�� ����{��c�-g�&*T�6Hyä>�$���0\^�v���p��ķ	$����$�"!O6���n��2]�'�W�ē+W�b�p��$Ձ��y�=)e�T�K���i�_v���m�l�eQn�^=kƜ,�� z�f��@8�v%H �E�sR+X�	g��!4����KȮz2��ӳ�qu��vs��[B��.����us!�������r�q����*yOdr���8��0�ds��_m2�RK��҆2l�*�����m+��G���zH�X�����ؚ����o��3��|���y���;�g����Y)I��D5/]n�����P�6�7�Uds6x��"[����@UVO��!n
ƙ��J��Tj�pjce�C�=�i�F�����q'��^�rF� �娩0i"T^�	/p7O α_�لg�j��KW����8�@1�b���kܚ4+@m���=����������wg����m�Q#��0��M��{�O��d���������q���nQ`9K�ʧ�9�`<��'e.�#����i+��m��!\�K.zn�.Lɔ�B%�z��6����1K�7.�l2)�ŧ>]�?��U	b��+�D ��G�8����*�&�g	�鿑��ѡ�ߐ�o$�w����$3����:4���U?Ɲ����Й����s�~m���a�畧』2I�.e��q~ �G��~�,�A������>�$���=Y�O�j���A_GZ��������8FSXx	&�m87C��mj�m�)�Ry���P�K6�y��M��[���`�t��w2�K���c������.ng@�N�qT�E�k.kZ����E�ѐt�Yn���������F���~����|�o?�����,��X�)��<o �Ch+]�H�3��������J��:�B�0�����W����0�,u�1�	㪗��� J8Pk}Ϫ%�ب���]�)�������`��Ō��@��B�zO6>�~�xW58�V��x2��_��n����ӯ����D^��؟:>���s鍼��N� �m�
>��
'���X	��X�#ɂ(zW��!�yP@��g�JVsZ3���ō��A�@lC�D�8�8c��:fxcb��5'��^�;Of�<��o�M�@�����d,Yi�,E%��>�7�V�~�M��ο���I��5,Ѯx�"%tgv`��Lu���B��8?~�r�@��댻�k֞�P��tɱs��W+})�s�ӻ���#�D���˂���@%��'�sZ)&�LL�w��ptL�͵.>~~�=|z�n��|�`2	x�}�;�& 	�;�H��a��,��&9h.)�i׷�no��DK�#ʲZ�<�������i�9��E��{6��}�N����3^q�#1��Ȃ.v��Q7%R4v�;�-�R#X���e�d���q��A�z3n8���t]��oikh{��l�}$���М�]_EdoD��7��h!��[ݷ�7|�.XWYlS�C�.��&����?�����U�b8yCÎxQ>7�m�Q�L�@R��?�(�"�m��k��2�;{�%��^�r~g
����$�8�\�ɋ'��q�M�o��VB��n��v��s� �<U�_��<��f�q�(��X�S�B2C�k��ʀV��b#o��1�
�s���j�CYKI� �/�����y���3�?G��z�=��"�}�ȟc.�|ǲ̛���~l�w��������a���w�j�_1��~a�e<�@�q ��ݹu_ �{����5GRb��f��&�������S����z�Y+@�������=�Y�����I���{z�4k\��8����h���;�2q����ܜa4d7}8�Ϙz����"���òӅ�/��\��ѧ���>��a2�ϫt����mX���4����jkk��ƃ/	�~�ZA /��3�2��S*#+��Q��~����&6q ���ȼ s�;'�<i������q���CX	%o��6c����3�����j=>{?iP�뼿�=j?����q�i��(5x`���>����}Lʇ}��l/�s���!Jo�ڌ�.{�������	���p����]+ f)���nh�cˈ�)�����wz�-e썊����&7<}x����I��nh���z�_wV�5�[3i����^�;��ĳ�@�*�~E�c3�U���N�n<��7�O�Oz�i�����Egk�ȏ_�w�7�z���o��������*��?~���T�A������<�T�t��><7C��Ir���eAC1��� �}����*`��qO�^�|3����O�As(��םM�:�kFU�/0��U��R����'�������:��Yw˼�!��^n��0��!̿F�^���
.��j]��e,3���T�0�D/s.�n�S�}ŉ�4C�v([eE�����������|�����5}^��<�\��vB�2�V�.��<��L���	� ��ӳϙN�XG)�R�#y�CV�M�;8�&���J���G P2��[<��i֝)�Ľ�r�����!Er��<=�խ��d�=���2��� `$̲��P�"�˵�-P(��QW�b�{פ?�e��:X���% f�������cK�"���wz]U��Ç�͡f�W�Q��M�o��l!m�`5Z��g��._�B�#�K�=��ж jW'�O�/u�1i����<'���Q\>��1d� ����"d�d�Q~G���?8�/MeB���uϮ���L+ xA��x,h�c293e0)�D�G��n��A@�hs��Z�ZE��,���  Ì�A��l�U��y�V���zm	�d���W��EdX%����O�v�-~4����i[@�J�+��ډ�r�J�R;Ȭ���B�.'�?�)f�9E�$)��L��rg�d�g���RSl�<�� ��9�����5�"��N��w�x����Q�^�t[�����G�"�J5��j�΃���S���Č���R�opI��m��Jdܖy�i���6GSMY��:�刧ѕ����]��V�⁅��6��*xG�	{��lĠ<mg������{���O�W�r?>���ߢ�Z
�|x�'�0��r,�IO�?@�0��6�������?jڗ�08ͅ;���X�	G��[S��E��¢�z$�ӽ����p��=V;}�o��s��'���Ul�82x��)�MVn�B��q����k��lqk�
���,��)�����<?L� d׆zp��U.�ĻՑ�ؽߴ�w]����j�l��|'m�!�ֽ_pT��I����/�ԩ��'&~�z��aw�;Qi�m%���,�/��<�{�0���Bॖ��XH�������[V�G݇΂(A7x���՘��_�!L7��.�p�`c��\��δe�]F`��8��i���9����`�Z��5���U���Jփ��s�b�ZH��"E����oX��ד�ɝ�����|�j����ׂGdRu��E��;Ά��DҸ��9�12�Y��ys�W��qn]��؟�r���]]��ԴWo%U0m��`�t�y	�7���o��Ֆ�=����=����WxS3��]*;6c�N�y$���J�+���H�s7�v�DV��ss�� �rH�31�u��E���P��@�uUKpsRu�ϰ�o��H3�}|�R����G���j>{�����aM�	�|e����:J+֞~ �'z�s,�V�%��`z��%'0�>!P� 
�����1s(�̍R��B���dk4�q]�^��|/T��7�eNJ�\Ż3����y�u�Y]���߆H~��^�
���|�7�z�Oҗh$���$�K	IvhWɚ�2T���y�{�]qH�z��F��PA@��5a3�&S���f�\�乀 d��,9�(�ދ��ʷ��ϗM�+�&Vu,��b�K@	wP^rK��}�񨼏�i��x<�KE:�t)e��Z�� ;��g�_��*�����R�Zom]�9Ŗ�s;��L����G�Jɇ�%�ߗ�}�g%��v�/wf�Fs���|�;�q�m�����f{�x��X �"	!y����ޖ�4a/d����b�*��tta{�CWn��(��`7T�~��~�Q�Kz�4���
�BJ�9 -��j�g��e!��B�鸏�؀�V���	�)%��]]	f��~�H+��=K��h]`Z��XF�Ȍ�)4ή�ST<���[\d1�!;�p�V�2'�I�����Ǡa�͟E��9�V`��\|H�Ōі�?b:N��K2K�<K&��rX���,\�2X�e �P�(�!d)��á�c�T.^�7��c��ã�B+��o��9�^C�]�������d;?�:CJ�4�PE� �R�4�~�՗N�YК�Z�)T��8'�q�wR� �j
�1�D��ܞ�?=�J�"�q\�J�E���s������e���kL��ʆ���P�~Ū1v�k҇,A�C<����p�{�{�[#麄,s��{�+>�n�PD�,3&�����0�ō�R$�5�����K�x��m|k��o�}�K�3n=:���W5;J����ۓ@w�7�J>�0f��O����@ˠ"{�ӡ5����L���&5�[� ��]' YaNԹ �ʇG.BHi�1!��Q">߽�bJ�^�zqȃ�I�n`�<���,�?kZ�=l�6/a��H	9S.��RE�D�UWSsd��-<2��� ��P���i���+Z��"��_a���"�������X֜�5I��*�]��w��^u������ʩ��ҽ�M�\S"�1&�SZ�G���A�*����n�P�pcis�ϓDO� ��.�2i���)%����Κ�HY��l�)���H���6�$MLB�C\���'`]� �=6�f:#_,ǘ�Tq�����I���m`��h2���P����_-{�@4�V&�
s�N�<UǼ>e�Z�M~HO�_�\��d�?��S����d�[9ʶ����N�W�J�0ykƩU�:�c7�$�M/8��5)��4F�+(��"A�@Tݹ�!aMN*�G��;����]*�dL�%_�.C����=Jذr���R,�E�=wjd��E}��Y5�UA��ZoXy16w2h�q1Y��B'��'����1B-!4w�yɃt�<2g\I��*���S�:�N��͸0o��ò�t�=UN�~���G��C�tJ�������TOD�yW1۬��o��oDB�L�F�L��-��"i��0 !%$#\����g'!l!q>�#V����]�V%�9f�>�=`u�c,bC��pӍ����-@�O��k�i.�q�_�YǤ�]|�7��Γ�$��7�_�fw�z]�=A4	�jK����	����{ж޴�ŗ18�`"_�8�LMaJX���/���W���z�KӢ������J{sW�����T���W��n*��/�PPd�t��Hv<�.J���P^�;u��%)�����GL��x�LC��|)�T[�K}]ӡ��pl���/��'b��ɪ�"�˻
��J�Mj���<,eK�Ye#ͥg�1�5�MS�+k�k[���n�*\(�E
=�h�NY����/�_`j�Z���wZ�29"3_�F�j����
�U�3Y*��*��[������?r�R�8�b�y(S��(�zG��c8d�*&�\k�ݞϓ-}��ӝ��(?���!?�A^R,��7��$%�Ө��?5(���I%�:f:�-�H�K�Ԕ�{>6ջ�ұ���C~�G��-�^�eU|���MB�+wjv��=o�����3g|���*�_��_��dOE��
��)�k���2IHp��q`�4WbA@8��lS�$�g�09��5��>:^1z�ɽ����v
���ZYi��hT"!��«�P��'`hRm���/�(%@I'��]c��}"�>ݯl������,.Qzkͣ!W����B U)§)���b�8��~6ek�CGX|��?k��r��!�TM�U.���������-yG$���J���Ka�ħ��:&�bҺ&�Shw;�����OY$���VM�\�r�g��PTl%v`����[qU��-B�L���h�-ȹ�bZڔ����Σ�@��mX��	*J�1离g�����Y�ஈe��i�`|r.Ҹ��iM>�~�Jf?m��=��� ���w�-T�n¤si'��'S�2*
��!~ͺ[/�3��� -�U�" g�i���4_
-��W�C_�i��������rS��STJ��U��'��	�U�sٙh��`��G;�Gg�c��Xȳ���g��0�/��9O%s$��~����-�o=E>|/s�X�G}Wv޲@� S`��Z�@e���<��>=��6�͖D�J�K|+��aױ�X��Z�����*�[������	�:r�TF�a�-�O N�U �8�|	8�L`e2�˦�N��me�LƳ���_T�����`T����w6����F��}�F���qe�Was�s���~~�h��1!D%Oh	1�[���|@��!ˡ���]�>��vO8�(���@=4�R�D0�)�����%��@�z���8��غ{nO��`_l>�x�4����I������|�:~�AE��J%�ȓ�YE"6)gl��M��f8����UvzM˕�	!]��%�B��a|��_.b+r�6�~!�3�p�K��0����~�+! �5]i�AKW�_�L<�N��fӿ��&���Yt���(�'S���eF�O^=�H7�l�)�:�V Wq�P�L�x��d�v���:��w4'�Wl���:�6SZ:W�o�����¢D�dT��y����	�<'H�%��d�D,o5�/
�N�������[��Ҕ^�dМc�q���R���ɼTV{�n�h-,�3r�Uq9Xxvq������6.�Xk�|N��g�ǿ�Hg�b�׌L\��E9�rf\�Z	�a���0Y�x
�e/)����(G�����?�n����|oǩ���W��F����_[� -6��Y��%X;N)�Q���8'r���e0��&
�T2��g���g	���O������O��!n��8s����*ݐ���I'�~kTc����䫁������Oj�h<cyc٧P�	�R�To$唀0z�������4(��έ�����9�ǅ�ҫ����낡)�Nu[��6�Ǘrh�� W�V1"����_gj���$,�^�6>��y��
eq�A������	�ʷ���Y�%�	L��۾�Iu=���BG:�?O��҉�����tޞT��a���I�cΊ���&�߭��a��s��i˱�n�Q��^Ryg��_���4dGe�\Khs��� `�A�F	��+4�;��5Ҿ���/Y��,�@^1����YxZ*���Z,)ƕs���~���Cۋ���k��]��A��#eKɗ��Io7M��hB(� 1�&�V&$�W��\���I4����~]^�9�H��p�TcT{3'�\o����a��ے�79����4�w�'���N������W�(�r-�ջ�U��S��B�90l��>3w��o}�r*J�8��3e��p/^�-BM[�{� �fu�p٣��j�ӊ%f��x�jZ1�C6$Z��)ܕ=`��ܒ����dVZE`�� f@���l�V-$?�F;� �Pl��s�B����f0� fA<rq���FH}U��WS�`�8��O~��A��Ð�e{�� kc��0��'�I»zn�Y}W��7L<���� #˘3`$�[?�,�B%|EHh�OI}$�Q?� �. ��JM L��bT���O���<M=������|�m��y��&�S�}I�%͔�62AFȨ2�Df_,@�YC?`�j��2l} �m�5z��T��JCj��������7���>��T��*����$Q��&�9iu{�Ń�K,���ڶׯ��f��
R�Jx��)����)/�!��8�P+�j7�#�� �]����P�<�ѥP���Nζ2$��cl�ؓ�:�DI�yAa\�I�	�++7"�U��Y�j o$�;�0��oû�S�ٳ���{$���r`|���A���۬��1����)��B�������wS1�NZ��M<�9��E~-�����P\X��sÌ=5q��w��7| �z�r+`�:[)��J��Av�����sb���-Fn��YY،��ʟ^���s�b�Ү��v�@�{�w���*@���F�%���'��*�6���Pg�\�eX��d���<R<t���Rg�O$mm7�f�ä��)���3m���h, �-9�u��Y�����4���8���|B���]� ��&������n���S;i�:W{1h*Š?y���ʔ�n�I}|�w+��b?�U��*��=`\���⃑fH
jࢅ�L`�0��A'��H��,�1|�t>2�S����1���J�%��e�3`��n�ny��'��8]̗W1�MI�R�8������'�������&��0/���lƴs�I@#c�2�{�~������	;��a�l[W�^��퇿�<	O���~��T��t�����$��PYXBj?v8mP!�K9��#�4��Ex,����/)���B�w�����5^lE���� �W�������%J�{� ���V�0���2������'��d{�gĔ�����VOڟ-�v<���Wd�ZB��A$Q'LwD��UWYo�#�f���q-4����$���
`�@��(���^X-u���2�~(p�������|� �����a=�����#�@M��=:!"�`T3���-�(/o�`ϩ)O"���_�곀%����E�v�4^�͹l�U΄elP��(���G�U=2������Y��?��r'Th�f8��РڂW����œ ƀ�j��h�e惥���'�����0�,|@U�A�˾7�|:��J5���"�!n� �q����  �9H+R��6	kMh���;�Qu3)� �$ڀ��Fʲ�J:ϯh0 ��	���>���%I���vv���F�y�P����pCO��XF��#m�\9�����}�@����+E�O��^�y`���q'}�̮�"R�C�dH͢SX��Я�+�Y��5M�Q��>��4��P�<0����F�s	bK�ѫlX�_`�0�c0�o!n��"���^�ѯ��ҷ&�-��nJ]��W��
+⯉�qG;7Ǆ27
�"c]���$�h��0�l0lES��>o�˿��)�������� �a��Q����:�cy��R���qU�R_��u/�����R�td��%��K�X`���I�m`�XR4J>�������27��E�qY��:��fK�=6��gR���P��	�Xq��v���Q�;��U$�.��'WI��-�<T��D=�H����5���Ks����)�!]@C�&ϕ`(��sc}��HR�S*����"��	:.��w�H��]��Ɣ&��[A�qE���,�!�9�d�D=��$���l�i���(#[�p��]�Xf���Mو� T�C�R�*Gؾᯄ1���(]�A��TIR���s ہ� ��II��v�{�x�YO�A?�l�U$3#�aʠ������=�#�����Џ_X�!���xj�#�R�2���N�=�N���2�P�w2����? 0�s���Ϸ/I��u�6�@��$	��F��0��Ru� N��Q���ʗ\�8���t������9x�ʽoqmc5�a��80���&�DOz_�G��λ�y`H="�!�D�#�q�H0J�0��V^��lr��0ln"@ 	md ���E%^G�G��O���u��3�O$�y~Ĺ	��p�D��ň�YU�F���\�j<G��<�0���zjuΖ	$ѣb,���x� ��:�"�䏄����y �S�Y"�����D�SF�	��J��)���O#���~!__�ƿ��`��0P�\Z��6cי�LaP���m@@�9�)�v����+D�-i>��
�11�L2֔dCANe �B���^A�DҊ��F�Es�h����V#����l�W=�h义�筡�$��g���Fd�!d(gPҵ	���{"���.hЃ�D�|�"�8-�P�yH�{W���_hV�Ƒ���Ͼ��1ܹw7,0�A�]E����ku� C+�IZ�S&O�{����͍����g�d���=|�*�:*��K0� NSe�&�/z��05m�DE�b���Ǭ���66�`�NE*��H0��'��b���v��� ��< c��ڈ^痑2Q�XG%����{����ً�ϐV~/0��`l5�! �s�# �Κj�X]���:��Er��!��/
l	``_��W�B��}���LA�BQ�Q�.8�B��F�<�d�Ihu��l0xN�Q���ؒt�ͻ~U[E�K� Y|�dQ�dKk8����$�`�k&T�pj�ȍF��;.#� c�����@��.���yT�Ӷ���@P&�X�"��VR���|��'��i��g�]�+v\���vߦ:���ð�p2�A ��l�Q	�ї��H�@��6K@�E����6xf[X��#�4�(u��K�B��^d�`��c`P�b�YKe^1��-�k/ѫ`�7zo�����Ê� r��;�
��3٢���n�C\M�`S�O�S�I���==o�:�V��'��;�?�`��c��$<�Ms���Vܴɕ%^H�T�.J�`�N�?��D��C���uU=����Ӎ�J�� C��G5M�/d������x0�^�5���#ɩ������_`D	� F\�y}�:���>E^� ��������_��y��t��W)��POy�l0$��7��ч��K�}��b�VX@���>�_ J}~���/���`�sk`��vq�c���-����'������NK����b�1][DE�R���4CvN��6Xy*�[`c����띺7��_�j<�t����7�7���?����Mu0. ��`�e�H�.�t�ǵ��H2.0�������y���zn��3� b1����}�D`���}o�.[V�㭠�k��M��xP�a�0l����=eOR�nZᥞ����}=V�L;L�lŬ#��c�iF�H1�[� �m��{���(��� f��E�ǹT%� ���u �pI��:~���Ϣ��N��v$٠���A��=�Jt��ZQ�����/�-V�``t0�^��-��F�$�X�+���T.���C�҈C�T0�0��N��J),0�ы����	Q��\�5 ����Ф�T���-v���DH0����b'ɍ����� \2$��0����_5��إ}�p�'ۓ�
`$F�5N��N��V޾v���^t1�7��NPW��ے��)�i #/�A�g�>�B`��c�:���t�D��>R\8�p���л=�� �fB�fC�N/M�%T%��pP�1�١�=���	}LR���������J���:Y.��� �G7�#ǵ�T$��a����o���D��LE";���ɍ<��ʨ�mI������$~���k���dTE"�|��o,޹{Ü��n��.} i�y���`�,P�=E�1������+����|YCgA� �N�1�u�����v ��Y�yJE�h,��\,b�)��N�����c��V�0��.&\�It��}=�=���JL��!C���-8��w�c�v�8��=�M�H��h�O 0d�Е2��I�=�<_��GV�r��������(�s=�ӂ��s���zN�)9k0��b��S��U7���m���<֮�� ����"��-�GLE��_�Z*��R�6��|M&���z;`����S*��$�u�\��W�/��j~8���1����Ǟ3r}�n����Q��zI��$��2|_������0�9�^ۡr���z���}�3vhq���:8�lee��P9V �� �h/��R����>�B��m˩���pS�n�=z��Eb߈�A}~u��z_������My�%R����;�}�I�@�m�}�"Y�ĸg�e��<%�C��mtn�������1մ7�F�z�=���K��0�O�$�XQ��)���q����"����Ͳ�HD��ɂ�k��Q�~���V�'n�t��N8l�;�3-zĒ���q	F�ȳ�-�
[4Wآi*�͵?�V��)��c��`[ �K��
ze�y��&\�%�sJ�U��tyҷy���w�	6z�d@�����6���S4�������`'ρ��l0ئ:�'�2qw���LҾ@���A|�:��e���S�<�:�s<S�6s<'w�8�t���u����ZW�ۀ�m Fw��
.��=y� ����~��M� xX;If�=yv' ���5�=��e��M�ł��y/=����z�i����7� �@)�t���
�����Xu���VG\ �����s�o�[:]�0LE� ��hN��' M�e���Z��,�9 �  W��a���������%�n*�� -^�{{{�Un�0�γ�Y��U�U.���s��W���<_T6E��`ȋ��y;���{9��R"��,����主���ߞs�ݝ�8�,Y92|�]@5�T�
��0��T7�P ��*��F�>�!��䩅��6U$2�lVNo䉷��$0ے쀲�sg=y���6ß$�h5��W�Z����V'�ܥ"�s"ŀ.������=�#1idL�I�r�_�u]���-+R� ��)�8�t�N��LS���ѯ�@+���"���'a��]�a<��lN8��?��}T.�=`��R��f`%�$"@�N����= ��$;�u�]�cG�l�_�;���j��O�)ʝ�v��8��?M�E@E��ݓgM�\M[�������9	#:�mB�0)DɄ$z�y��$6���dؖC'�t��t�j!�d�_ ^Hp�.��+^ٓDCF�թ��:yU��8�#�
g����e� ���=!�@����3��Иœg���q�[g|���\`R.$�s�K0^=4����#q	�ܗ0�#[�`�}��nU�	�m��4�*f��I��!�p�B̄yQ�F���0���k:��n�m�m��c�݁i���w�\8�x�H.��2��H8��)���;�;����w�Y���9ڊ��?��m0�8��&|�ǳH0�|_#�h��F�:Mj�%IeR~�#�w��!"�ci�g���'ftЙ☜��Vl�*[I3��`�\����2H���Vr������"�,�)��!/�:��^�WƩK1^Ĉ��m����}e�r΢������^{�8�{|Gj���o5��wX���JE6�/ru-pu}��L�O��k��}y��T�h���CYuM>uъk�\C+�����]; ��4�u���|������
䤺Re�*P7ĝi���X\1�ܕ�g{�Ql
���Qm[�X�>��w���6'�gu2"З�w<�c�t�Z�g��#r�0_Z�m5�%��yd~1��-����[�#+��F�XW��S6;+-O��hK�3`����9���;\mAQ����]C] ����1��tO�ӣ��"y#٩`��4G[�֗	0�70>�. �<�6UmW��V��
�'0��<W��-������l�\�$��H/._�b'�^������E+�Rc�XG��9A�#۟<y�޹�ܽk�Î�WY��u�5�C#�����\�A���n�O��Y�`�����,�����00�P;�Dࢩ#�:	��F��
wO�xm3O�	A2U�)�uZg'��o���'�!��d@�(�E,���t��A�E�4�,���uY1�9�[�Ic/�գ
��,8nɌ�cҕ%	�p=\�&/�s�[ �#�K��No]�^>ˏo˛�}}�i'���WK�����������i�Z�:�=��gTy�x���7���D��@J�� CD�+��,QB�/�a�D&����e� F�C��`P�V}�?`��TE[����a�E(�X�A�7�����qXp�(LG����/@�(�mV��h�/��,)�����A��I>J/��i�$��ޖ�x�<�!:5��-�e�8�t�=�'Oі���s^�e�Y����v�qJO� �<1�ԑ����x�s3��H��.��0����p��M���'<���ܖ-F��a,U	�D� ��:��֭[��-�vV5�#cc"�im�_�Ԉ��ה���<+U	D��N8���D_���pq��y�'OPk}K:0NV5#O�(��<���H.\���e �k�G�!��\rHI�S�2 ��8&�#GT�� ��p%}��tmEj�!}��߰��8w��Jp�@{��ֳP�-FY_�}j��,�V ��h��d��8����`L ��T���ƨ7�����_���[�:1g����kaxf>�(��Y���`�;-��!�_�j�+G�����a<�e�I�]z�UeC� ��	���L>�~F��#�E�/��o��`[�����h�T���:x�ʷ�ߵw⤗�˰�.G�M�<�a*�h䉫�֢���W����E���Nz�.�h��F��Y$��<��&O�V�s��Ƴ����B�$�����3�H�.��A͗|�Q�;C(LMM�h�B�ꫯ�ME�xBo�bgA�
eB �O���zDE����������]g��s���|p؍�&ƣ��m��s���,"at@z��<'�\�Y$�"I��m69��q��f����C|��盬�db��*B��1��+D����%�O�"�4�i�E���ޞ<mK�<y����)O���qR���&M-\��$�¦E-�x����w���D������.�"Oh�M����T��#ң�L����0zQ��)�@j�y\``�>�v�>
��6���#�	&.6l~l{�.�䑾Q��8ݸ���ek�/u���%�ψ@���\:����	BW�t���Vކ�g����a��ðî��5k*�ߣx��w�K@�-�c:N_���Ä�*�H��6g��9�v�K��g�'��h�v{�����
/��3�`xaz��Oy��3����ՓgR� @��9dr>�
�OfЙHۈ8Bˌ<O��30��_vN�$�#hS~Tspz�Eu^�z�o2�'R�w�M��ٳ@D�1'�JNF�v��2�j������?��o���k��0(�����1֠ԡH3��hUF�2���P<?��9�4�yf����%N�8.�Cb)m�Ln�<O�$�D���	l2�ɕ{&~s/N�P5ahXůV=�r�l���:;�1��2�L��"�],�Z(����/h��'uD��Ǚ,^���i��O��`�"Y��'�[{�x��5���%z�zG_�L<|��>P�W�ԗ�����
������S��c4��$g/��FT��4c/��X}�@��.�(
d4 j���TD�~&IG�~k�����Q�|:o7�|���'c�24�^��.L\�VB�I�|��	t>s	���J�6�O���[ #ߎ���v���g��s?:#�Fq��� }L۬}y	��*Z��I�r �S��������_�vN'�^�7�uu.�3����zx���I&�!���K��:��tի�u�7R
={��yh�7�=��$�E/_����$�g�,�m���W=�W�_ck���I��( �Xǵ#����h���%N3��`�;��k���3���`0!S ��9g�.����1q�u�J��c�aXDi�Ő���J�1L+�$%�c߰�;2*2����Z��Y�����Y$흛�-���\mY{�DF��Ú ��ғ�/�_Xx�W�k���S�QY�~���Xx�WN������sY�kI<V�X}�K�q-��/�����`���X����x�\Ց��G`�gGvC�T�J�L^1���I�i?�A�~O�'���3�ᧅH^�/��ʲw��k��7_��]:g>HuB_�N �oY�����<��V��P������=y��m0��3>0��l0l���?�k��I`��-�<k�ń-�]%195i�.n,��~�m�)�l.P� *����p��m�0 @�򷯿6	��b]c�5��0���0�G�������0!�z#Z�^��$
��~�V�˘W<��i�#�r����T{ǵ�)����p��p#�����ɳ��,���m���?�O���J9�}�X;l'�Y .X@�͚�,~�w��U��a�D�> ���>y�!pQ[����+|B���(�ꋂ����@ ,�Ȁ��s̀Y��9����+p�Tr C;HF瓑�>M\��t�T�r	^6���%�@��.��go�$��lO z�x�	�� ��+!�:��ŉ��g"�ŉ��+UI�Ư~eq`t6`�j��N	.bED�H
�"��
/���|�#���K���<y��w�he9�����yz_g|pV Ck`��]^Mvy{ڮʎ*xcF��ft�: ��~4����ѣ�����R{,-a��$���w�}���D�+/_	`H=���� 6���ɓ�w�����,����B�<}lj���_���]i�r�>�j�K��s� 㯬"��n����<9�L~0�*9@j�l�8�NIǵ#��`�r4o�Bq�X�*��O�4�u�ߗ��7�q�1 FT��]+r6%_"�$�"�W�Ф��~l�&E��0	F%��b��z
��qZAF��ȼx���<��4��RQi�{8L.�F2��N��i7�L�HT/v��}�+yR^0��$0jFIq$���Ĳv��$�pФJX�["���]L�9ݸft� 
��$H�v&�H�{�����肤]�@F�g��?�U�:]�:Be�x�'Ok? Ki�ӕz�-���"�<y�������#6/Ο�V����~tV;�  @ IDATj��*��{�H���0���V`X�C��HsV�0� �:`������?��/�!�I
���߅o��V��&�����(������ ��?��C�A�Q�*���	㒎 ^�gƓ��`����(��4:TE����`�jF�qDpg" ����ǔ@>	��p��I���a@2��<=����<ߣ��r���^>�����7[b������e��F�� �8�<�"���wM=����JE�XTS����ڞ�gi==7x�@�7�=�7����2��B;���>�(�H��OP>����*iZ`4V����3^ Z`qܶ���e��F���``dk����ad�����Ht�����L��@C��gޓ'�ƅ���gQ��������g˓�=�i���!yx�������׆�2�l�k`�����%3؜����C���7����x�w�^�׿�e�!nS�2� �w�aW�"���� H4������O?ZZ����B|���Ev�`@�������+�!�� ,r9�D[k�	�)%�ɸ������}���F6�k��o�G~���� �?ǰ��X�-��6�<�������=�����8�Ѓ��k��~��uu���ډ�`dT;%�b������0� y)�6U�<״Mu�ţP�44�ڦ��IM"Zؑ�E�X�}�}R���v�PA�`,,J��h;��p���e���@^'
�햗~wߦ�~�jV��
<<1�w��(���MZ~=���{�h��T�T	��kFWQ-����s�Y$�8��!@�ܱ�#8\�]$�R��"�m��R�,..f�r��������T$�[��i ��7)ƕ+-�q���ǟ�Y!?���茻q �C�%"�x"u	;Th��@��T��N7hƳ��d��h+O$~k�P�z80����"��� ���`�ID���:��o0~%g�������=O��G�3�+��ȦN��_6.�pG[U�fh���Ueb}>�����Ό<�0��)�L�1ԯ�z�̈́�����W���˿�
P�H�U��u�ɸ�`��'6��Sj:+���
�H@p#OmQ]}���� _$.��_�-z����Y*֝-	FS���m4~?��P�)�Ѵ�Dj6�rli�h�ᓬ�jGjJ��Vޓ�ҁ��k_A�Ot��Uj� ��y����V���֗h��ٯ���{2�}�NS�q���ǵ÷r0G���r���U=�0�߉v��yQ�20�O ���'��kGɆ�*��&?��C�^vW�E��@��m0���_~V�E�+ڮ*�1U$ �(�x�8��<��� ��\��0/)��*\=x��� ��cx�"G�6�d-������'����Z蓛�{�b���v��:���uN̖8���L}�К�=m>�t��۔m���=�5�'�����	#V0" �\@�����|�M�������h޷U�W_���~�3:��t�h�T.�C�B#��,���s��� ��`���WY\���d���۔�9��.$��{E�O�:CLW�c��OZ��l��D'�~/��Y�挳1�G^��H<i�1;��>`�nJ�4��w��n�(��?���׼�04V>9W�iI'�hp\������-��#1���(Z��G��N���^����e������n�<"�o� #�~��D�:����qN�ۿ�[u�_�y�8�	X.��/`ء���I0T8�b�`�l�0���W����:,pC6/0~?�h���o�.����w�Ib�H�s��Q�?��� ��0=5m$f�a*�"�Z�i�2�B�B��y��8�d,'�a���$�I*�<��7���.�3� 7�};�2�Ѽ{��ķ�tNX�����%yۘd��Iՙ�:ӵ�ā�9I��x���L�@xN]�0Y<\E�?*O���1{�<Tk��ܔì�v�Y���բêT��6ջ�,�8[E��6O��3Ѹ������e���4��Q��*|��F�g�"ɵ�jI��Sj����a��ݰ��Nm.����7uPY���Y�nǧ�E:@w&j���YtZ��W�D�����|��I
f��n�8�?V�ڐ�E��䍌��ag�%9�6:��-*;�+���\���ٸ���q����[���Te}r��I�.#��Ʋ��/��>ǵ�R����8��D�ܥs~�92�Y�㔡�0~���k���I�ص�O��^�'O�e��$k�^���sH�v �[�ן5�Qc��v(o���6|&G[Z�w�u���sBr�` �H0"����������$ �Һ�8NS�Ҏ?��3����'�H~��'s̅�-ܑ�F��ā�q:F�ƿ�*�/Ǔ''�0J�����VJ00���쐅;~0�p�2c ��(�%�(\T$d�ʐ���j�fn����'��"�����E�]�.g�������$/�b���~��Ս<��i0uM�j�E�/u��u����E���r_~�����v���DQ����R%�o"Sۋ�{V���bQq�egLM��b��mW���|����˰����ݰ����_�|�+CWNCeѰ���V��]h �;�/���AV[|�10;i`�=yF��_N]���N�\;��<k:F�!5��7+yh�%�y��$�<�]j�4V���j6�-�����k��/���� �����I�����]4?�c���w����zZ�>�X�vP��_���{�g�����_OY`�12%��l��6p�q�@a� �t�p�`����T�O;+�ˡ��{���&�M��;0�u ��O6lS-n乫�^���<������Le�#@�����4�A����1�HCM�i��<�����ϙ`���3�� ���B���؇]����u?iv5�F1�I0.prT���Ȑ��yL	�k:�Ow���ք%?��)�|'Q������B��	�Q��a����:ߚ�X��y��]K~�����F�xB�a�9n�/S�`\�̹��K�' �P���r�$wd�B � ���&^�d8H�\?�z#QN�N_Bv����N�i�U��C�1"��'��6Տ ��|�,l�~f�.8��qal��|{c��_�'�Uݸ0��"�QE�1�q�K�ꇃ��쏾��o^q�Q,�x�-�Z@1t���O���(��ǻ^��������h�������p�֯��OZ���I0�4U����`��V���x!�5b�S+�r�A��Wb���<��2bg��T�3�u��y�]��I0��0��(k��0�ǔ`h=�K�ѧ0��:/��g� 0�bf��cV~0"���mE���M�_ڦ�o���հ����~��v�\�6U���IB	���3�H1���T'���믿�_ME"�Q�`<xp?<��H{����@C��;�$>g0.ȏǜ�����/��q�q����B�":����x��5���'g�ȸlOGh�V���R�S孍Ú�4ihWS�n6e�є�"|p�qC~0$'뚍�c��I�pZ�yV*�!�а���c{�4���̤��LlNSKx�r�އ�`���%����C�ʧ��N�����r>9��&>��T��G�d�(�v��m�E��95[D2��$�C�sLg����4�_=��k
Oz��.z�&w�x��3y;��o��i�qO�<��m������A:t��+�n�Ѡ����q�:`�N�іhc #�ϸ���gu����	0Z6�I�����@�>v0�;.�;ֻ��.��oY%��c��O����9�G@�Ɗx���3��QR�s9`��Z��D��lw�{[Y%"��f4��BM��Y��H��'����S@;��1���GQ�,��r
��ϥ�"�Ome(�X�x��-�M���f �O �,m=ԛ^[�,
,Ԭ�e��~}��D??Mu_�)ܓ��̴|SLg �h����M��r�����T*.�h���h�FX�q�` ��]v�Ƽ�����������sN�^�\���;�"'�;�:��1W���$�4~��GI���O���ȼE�V|/���V<v[<b_k}:�%�
�4�=w�V�BM�ޔ8[��X6c@�p���R�E�"��!�6Q"��w\�����G��0`$���SC�E)�gq�������Ƨ1k�][��Ky�)&8�9Z���-�x��)0p��c�G�ئ:1c��\�?����?�?4ܾHKR<����%��[~&_2p��H��Ǥ�h�M��(��I�s��#�A��gϹ�q%���2��/�VU�H&��L�˦B��lSU�_�wV��Y$�G�� �wd���Go����jрf�����/�?�j�+D0�M��k�8 �1�E�Y$� �)K�g��es쟩_���1��6��Yח���&�Y$u$0b:�N�l7u"_�� ��t1���h3t���`6��{j�K��jg?@S c��7F�Aql���� ��ֹ�����h�K���OR���k�E�4F����c�o뮦!Ɔ�D+�4��s4�H��[\�F2�͍C2Ic�~�~��P�\�|�5��:oZ��gq��M���q�vy�u5�'1!e���}mF�ڪ�/��_�	}5y��d`乓��9��xsQ�-�_��)��i�6�u����TKo���믿1��7n���6�`����3H0�x�?U3����ǐ���s���pW��^���F���ؿ�@�|3�1#	̅�_#���U$ƴ�˭���+�4�[*��A1[��j�A3v&�z_5�%��	��ݨ�=��w}�Ӑ[i&I��~vO����S!ɐ1TS�$��F��oJ��N���Ĥ'�6�&J9t�g�xǞ!���>L���p{z��S=	�h�߳7��w��ܳ����lk�����/|`��c��Wt�U�����%��eՖ_�������ʅfXƯ�~b��T$��<ݩ��р]��~�Ri$���G�D3���&��'�8��\��=��X�/��b�)�+e�0�$cR���8�-�V�؇�E�Dr��v7V�pH5����i�~������1�I#�6��}��mh�h|�����x�� M��h�A>6�iL��[''�ȹبv���A=ҧ��6��"!9�c��S]��u~�yB�u�K�x%W�2^�˾ .���ƨ�����c�T/[<���%N����B��OD��7���uR,K���+�z����e�4"�� x�`���g������4a�Zw�ޅ��Wak�u�m���b��n��'�O��:Y���f쭪����Z;|�3:��%���C�3�)��%�E����ڊ>�O��8T:�b��sW����<�w��L����s�=�Ke�6��ĭ̉|LXk� FUq��c@�w{�����x����#D��$�q�F��wO⻕wr�%U�$qr���ή]����aQ�Y�^��W/_�[�
޺67�\K���߄o�іp���8�{���+��R�,��V��w%�o ���V�3"k煹�"�9I0�.d�1��{a�=�Et��Ŧ���Z��p��8x�i�"�a�����<"�5.�W�z�Q������W�&�~��Fb��~�>잌;9DJ�/,�X�{03���\1�9�k�+���4�l�2d�uW�ڻz]�������N�tJ���{��4���)OgDS���'��b��L�p�5��t��vח2^˛�+�����b�-����m�����~��D[�MN<c���K�|*�1r_hd44�Y�C�g�a�,15�{��6�������}�j7��N74���jA��|��>���݃L�)x�3`�O��yzޘ߾P-��Ay���,;�K��3���.���Nr�z���h�*ِ4kC�ߓ�b_���S{Yi�*�չ�Y-�E_�M>4��	]�����.I��2����ʇ�P���ѱ��T��*{�,��wi�e��|��u� A�Z�Z~�uT����vBԥ��m��=�mm�X��#���o6� )�-Ҍ����ė���������\K]{Οj��vԻ�J��,ʑ�O�3�������U_�	��`6wÈ�@Ǝ\�c�WN�GGM������tp�SR�p�*��/t;F��%�@}� ���z�Ƣ�ѣd*�mݹs�"y��NLL�	��Ҋ�B޼�������S(X ��9C�
�a}:��|��J����������r�/I�A��|#�wr�5(V1Z�R����xdL�v4�ZܪW�F}@R���+���;4�:WcN}�VK�"�j!��KM�]��'��1W��9u1�ք�b���:ΞQw�g��}�
sۻ-�N�4��~�D�w��i��K�6�-]�����Ą��L�(KS0#(I*�g0��$M�X^���&�VR��^#������֚�հ��N_i��jI�����r���<pO=󡿼?�/����}����/W�b���F��l�CIƯ��ߏFV�!��Y�5��_
��Ə"Ɖ?�K��Ԏ�����z�yZf����m$>w>�jŐ�g �ö1SNR-x���J?)��ҫK���t�  .�E���+��.��8�=��N��㢃�|�xI�}�h�TG��F��_�G��y���:^�L��6�`~<�$�X_(|��ņ����̅�7��4j�~S�����>�"�7�O�q(����8<V~�C���~�.s.sW�`0o�뒑G<��m^Џx[��*��s�tښ�6�Ԥ�ɸs���5(o�R���v�` .��20�q[V��7��E�VD�eT\m�4:x�� �݇��!����݃�Bp	ܝ�-�C��.��ͻι��k��������~�+@�۷o�2W&��a�Y���^O>����c5e�ّ�@-���:�Z���V��x�񬏾�j�HN�2SA�	���o�yR��;�C�V�m�ڞHn����n%�!�a�N<Aٟ}<��Q��E8��Z� 3_c&�X8w%wI�|���n�iɹ)W�<	��"q�X6E�����"�v�\�bh^hEDik�7�B�Ƹ�X�h!���nk�K�l�gB��kj����??�kRC�[���H2
tdR#���Hױ]6yN�D�G�m�(p9ߵL'y���[��N���(�#:��٭gZd
�9L]#���G���%fٻ9fK�G�9pu[�o��B�W�xIB�|we�{҅���;VY2T\���c�hD�;Ӈ�ܹX��ο+��R����=���Z�gq��C5������=�5E��O�1�u[9dt�A[~ty&~ajh����R4b��r��p��~�aN���"}\߫+��\�I��1��Hx���k4r��=��2ZM���Q��M�8`�:��4�J�O��έ��.O��<DJF���U(B�x̰�*
��6^�v?���quR���O��P@�95EA�0`��2�{������0��N�vsE��|\�ݪm���ޕApW$3h���~���P���rID�D��j۶)H��U�e0��&;^���i��S�4�,q�D*��ͫ0��:�9.�(]7]*ר���g���Z`�Z����+��l�=�5����(������w�T�*���S�[�a�(�^'��:��d*j�L(&��$%�}���O�#�]���G�A��/�h���ඇ�?k��0>�N���e�	��$e� p��$�MtĐ�I47vzK>R����C�-��	�(�{%�2�f]�I4�"S�G�)��QK�fK���<��v�_)1u(�x7�?S�@f�J�r��c�jx��/}���A�4��*�� 9*��Y���Ϡ��{$��.�}_dt�'ơ�K'����g)����1"']����5\k�$Ж�/�>~̃S΅�ɪ���(�P���С�����&i@���4!ST�������ٰ)-3gE֝=�7[c���Y���?)���/Sf%���c�@��[�����.��_�2.YId(�1\�vA5ת�[�"�Jh�[�^�W��Sx\�P� .S���i��.� ��hNQ�Z�w|1~�]������%'��q��r��0:��٧�Qp��6�_$'7�A?1����w�r�-��ٜ�߯��V�r}\��v�)W�36�����R
:D���)�`�>x������w�Y(�]�#�7��i�2���R~[��a����/�k��#Er�b|5^�k<S:���Ƃvz�?1-}[J?��Cn��e�z�8^��.ԝ� �h䵗����G�P�1 �*t���>� ����)�i�A&�'�Bԓ,�dq���"�瀪5�%�M�큘��i4�N��>�U�,	H~�K����j6�J��zP��[ؔM�zۛ����ڬhz�|��H��V������"2��$TD�}�Ě�������nY5����ֱ��KR�!�؇��)2]���y@ݸ!Κ�^�zS#?��'}�������c�W�2P�:Pc״�X�4w�1�sue����M��2G�X`c�[�pFk���*�eL9[��t�o��wo1ef8Z֢��7�Nt�yn�����/����� ��M`�窂����Q/U�?�"��;���Ez��~_�wRw�~���]�BՉ�{�p~��g���-�]��ɶ�]�]H�؋��p�:n��1���4[���ˮ���#wz��_/�0  ���Չr��Q�=I���[m�A��C��~frQ7�"̆�ė9Y����v���8!Q�o����@��UG2X�X�*{O��9n��I3�<���e}}3+��w8n���{QExO�	�䒿�˩���B g�)O��*�͋kE���ᜥ�[�y�¥Ђ"�l�mW�us�>��^r��$������l��m��p&���OѴ��r���{�����olo�B��?O�Ӈ��S��*S��<����z�m�W���vF�u��$�w�ŭ�I:+}=�uTU_�/
��M=Z+�m�Cm<�o��:�W�mH�&���� ����M �7XA�hI,҇T�+(5�����Sg8��5$_1�­���P�a�$]�8smZz��`��\�]f{ U�5��Iy�DvI�^5�S�̏E	��~ׁ���!�o�:Il$^�09>*6��wT��{��v����գoϛH����V������h�\F5ӰK%!��O&�Ⱦ��]Ӓ@Χ|g� �>A�$~ïQ}Z{�r���s�������_cf��4T�L�gW~*<�YΙ�L�9{��y���Z�<���LxR�js��;��r;�����ݵX�ȴ��L��O���x�z��h�=%zp�]8��������'o
Ǹ��G�ߚ�վ��5�v+�� f�X�D�Fp��&o,W�y�-%���Y�e�:��ӟ�f��mY`�D��H�̉��5��<Dv�+�C<�e���qBC8MI��_ �e��>G��Usq���?�i��2�R�����Ir���z�hW�M�Y�b�K���k�.���%����x���6�y����,�܁��v���2L�%����Ë,}V���M3')4�0�+c�ܥՔ���`>�AC}���ֈ2�n��ԭ�Wdt����x"���s����e����$�ּ�����gY�Bտ3�x�c�y)� ��� �r���Z���� ���'�E��fX����ǆ�� �>�����W� &d�y�7*{9�b��V�������}�e�ɐ|�T7c�Ō\�S����9�k�Q��&ƛ��Q!,
R�3|ԯ6�Xnmz���ۓ�3�(�#1�A�ޏ�P��6����8���˲�Ŋ��Sl���kQgEay`���l�
�+�l��P���ve��0�C�v2zv^�2}�_���{HFj��9������{�Y�������f�ga��(v���ם�����Pn��D��dr��3|���	��=z�֐��f��LC��Z��=|b-��P2�&#2��������Թ	JF�";�x�O���U����9���B�>,��m�����R7]�.R*G䮵@ ��lJ�c������Ė�Y�����SX�@�Q�G��\�a��C��<XP���M��SG�1f5m�W�;� L�����Wa�hH 
 ���G둡'QR�����<��x�$���) ���c�'s"3b%��7���Y�x�h���˵�F�V5h�>����Y�Q�o]��������$z
��0�@�Rg�(������P��=x�m�h���"RK��V��~��3�X�^,�t�;�5oG	d�z���w�.�0+VYH�ʻ��]�/l��e�l�����\�L0{(<����� ���b��Geqz]����3���^ܐ�AE��S#|��=�(dB1�ſM���e �sq��M��*�23���-��l_&�o���o�����B�?'�&ŝK^��)�[6���i��D��~"^�]e��� �c^>�B��Ճ ����}�j�ӭf�*�����('�YI�ȉ��2�����Qu!e�#���������!����DE��<mʱ�	J����!ʢ��Yr.�+kZZ@��D5����d�Á?[��z�n��.��~�j�Q�P^�4:��4ÞN�cZ�d��'��#o�|P.��̯��$|�E�"�3�?D��QV��ܨ����b�m�;Gc���4�ɦ@2��9ES�dOU�-震��6��6�λ�����jj>ʆ��E��.�do+�U���&���������2GBp�%\���,����K�`3>�B�弪f��}M2Ύԓ	B5S��̆��z�YxU�Β���q�8�WX��I5�|z5��\L��$n���3����v�����Q>���3?��!�3��g�ٰ��,#Ɋ��{���{/8̳#�d�(��\|�	ہ�o$I�	g�V:��bg�-�Z��§	��҆8��	�-i`CG���q� ws����
����f9;3���}DR	�%e@Kߕ,��0�A�����E-m�sl)��l��a�S8��N��\�$�OH��>��7���0��3�
��;)��;~�ԲP�EF_bE�#�i>KP-�؁o��DiUcߞ^�=i�|������l�t����$ձѾ����ޅw�/]Mf*(tX �7�P�'��������p�䑝�$ ���ʗ �k���!��k�7Q�4�ۥ$��5Z�j#�[1����&|�U���E)s���2rq�6l�!��$��d�psG���pU�H�q��n�H��;�>��+�bo�J9�Rx�G�Ǝ����	<�/�:OL��E�H��8P���A~?@��_����aP�=$;8LKW��%Ȅ	E���?����]3ˋ@|=���<�<jFs'8 (�Y�_���[/��ڑZ�9�
i���#�z}$�r����1V@
Ƀ���~0H4ӛ���� 37����o�E`Ҍ��mt�.�n��G���R+Kd��_L�z�RկT����`Y�p�O�����v -<�X{�H`���+ŉaWe�[�]d��f�����H�7���!T��.��{o���䳉�((�Ąx)�x���O�L�ދ�?�f䡌�{>,��yw<����;8؛�_f���)�)o����̛�w&�nHv��ͨ��;﫽�"�x�@�~��%~D�wX�>&?���_	��K�s_��! ���h~��ԍ�v�!	.�OX�殹��&S��"[���zC)�
��.����ח镂ɑ���x�M�k��� 5l�4_��C��>5��k��2�!u�9K�î��3��\�]&c��@�$i��-O���~m���Tm�N��r�zq�m���`G[j����u��q�ho������ס\��B@��g��w��'��]�:��M�ţ���,?���c/C~ǣ��#L�,f_�U����9t;5��_�Ȅ����RO:\m�:G&YaC�gY��U�z(��v�������1O��[��a-M���^���~u1M�ZR?���,����i����E�V����<_���_��?�Uu�^�?��u�ъ�V�����G74h���e\�i1�X�;;ֿ����Ԓ��Kn-�)���x?e"NXp&(��^VI\�
p��=C�}��"9�%��N���J6������N�����D�贒�����;�~��-��:��(�)�R/��Ԥ��^�Q Pm�V�o�m�o�-o�]Ё싒��M�ۗ/t:����Wxtc���H+Q.GRJ�'��54ݴA��\��T�mJ�f�����$�͜�BPt�hPe�K�`c
�:��Ւ:�\�� ��?��O�R��87��/�t�a��	5{$�#��z�C� L��Y~(��Y������#�3D;�n<"�,,"���r�D�w�T�1!�G�(�L�n�BȽ�)jH.	��kD݈������KL�a;Q�q��
ZI �D�P�l���Lc5
���[3�U�G�U�1��6(���$��c�5�gL���Hg��A�������r#pO��l���W�)�U��P+wx���i�� @�-{���(|�cB��0�\�&I�x@i�`cc[A�n"Hh�Iʲ�����X|e�b�3����Zqbt�&/;|���S��$?UjC* �H�\B�މ
[leG��P+��w�-�g��ID�|������2pˡA:��$�N;wa����#b����s? �s���X��Y���B�����+�;�(�$iab�?��[���^�E����+�u,�V�3y�I�+��d���G���s���z7��m����ڣjb7�[t��dhX���t���Srh��?��qsT�B��.y��̶�b�_�P�����'K���m��$�R;���A��`�csc
�������=��n<6�6{}u8��>�ޏ8��/�rM1��9I��g#���7�b�w�Gy��k���q5ه1�d$��*����@W)�A���F8'�^W3��1ꉩ���b������c1�qF��ϲ�8TJxlVt�����_�6<�r}̹�t�$|��G$�p���#g�S����D"Jߩ=�N��|xn��+�s�8�O���fLSb.�M={�N��g����ä���z�M��C�����z�����Ϩ�S��DVn�eqS�(�fY���I��<䋆oI�~�[��n��gL�磻v�2�CJz\ǎA�R�	����diӎ�>֦�2�w�Z���UxL��>���G����{Ih�դ�ﯧA�տ�9ߣ��v�����>+��u�0��BݖH21�M6��%'$-e~�tP	�v�Pmf51
\�+,:������/,�]�Gو>�R���yp1���_%�^u�����}���F��e����&�ZfPg�ou���U�Z){�����Ge�ɍz�c���]�]�\\�qzX�"�q�P\Ǆ���u}s؆�Y���=M��^'���&s3�;'^*2N�L<sOM����l��9U�qǱ�kP0�@u] b��'��ď@(��<_���>y,�B汣��e�Ed=J�$�,�Z���Qs�A�E��}��j��)��4<C�Nï��EDp�0�)MR~	�m�|؈5��t�T&�U}V�$�6�_�T��
��6�·��mu�{��~��[|P�� ө�8O�=���b�8��p���������i�k�QR4^���S��*`Z9���H�IP�lCNN�5f�{��kƐ���y$��j2����ַD�#��`���F�1���;�R������aƉ��!W�a	1;ɀ>$�$!�|W�%�����%���)5<.K+��X��J����zt����9?V]4����>��gvJ˻���X�n�s��=�*�-Z���b�����U[�����L~����C����̯�+g[~U�a8������T��*g�,Yo��7�{�0���ո��.��d��S��:�r�l��܏YJ5.��쌡}�� Jl��Ⱦ�Z*vG���[�tp�|_�K*�]r$x��W�
9ȫa�����m��okƑ&^Q��lO�3,Im��	�X;1N
;�����TG����n�=���%��3%F$���gӴ�Bq1Db�j��4T��.�5ܑ '��0$,q��4ʋ�|���	vw��<���;O��5��c\��k�ʼ��&��>c��w���2�����QV�H�6z;�������8�{�Ǝ��b�v`��(N���/ׅ�>�?|{A�|�)��ތsG̗��(���q\!�x0s��-\kх3t�v��u<�	NPn*nn�Un���1��\I�(4�_�/?�o��|}|����{B�+<���D�F�����^ʺO�2�F�C�[����Q�lyp!0¬���v��WŕS�X��G����"�sVo�w ���wӆe�>&��b��ʧ �Q�|����)�c2H�Uc���M�.�"್�vq f���Y�1��2��z�{��, �Eh�b���b��H�պ��l��܎d����l o[��N�*9𗯄�/ʛw%�e��.Q+�wly$�kw����u��D@���)Q��_��LM�"'*wݲ��b؏}W�[�?��g
q��|\�g��C�A!I~0'J1��x�	���3��#���P��Ԩ��� N������3x�,c��n��=�C��l擢�V6^W��_��(p�� �������D��V���qiI*����;Qucp�}䌠�%VM�e�é��UOT���7���1|œ~W�-�}u�׮G�i����[7c�D�� ��C칦�A�N���(*��S�
�yC\�ґ뫙@Ps����8 ���G�fe���R��ә�kM�1ڟ0A(�����	�\8�Qx&?#��h=y�|D���t����2k���P'\�������"j[�88�2�[�ަ��)M<��C�xx�� ˅{��?\�ԔsY�Q��{���h|,���6>���Y��(и)h_;z`�P�:�l�(�nf�-��t����J�-�$<�j��
�Yi�wVr�i���;W˩K�s�S���d�Um�&}<P�*�P����otoq�i��dn�����D�]�BM�̄O"1HH�Z�n��'2���>r�!Y��R�'�#6�/�U��_��n�B�%me��1;w��<Ʊs*�S.�4:P����P;b-,$6m/��z��`W���0Å'
R.
����GǨV$�A�a����6���8E�Lw��}��L�����7������g�J
���n��:r:�4ӵt�=��jc]�@Ւ,�֢�u�di5��:5����[�E�@	@a+I9<�����x̓�}p��sӸ`����j�ވN�}��VvE�# �@�yӴD���A��� ��M����]I����Yk�d��d�(�!�GF���j)�W�HMV]"0�?�zC����&Y��M/��
$��V�"}%K�jjj*<n�.�*�1���Ve'Ue/JE7�d��Qs9:��g�m�2��.�;`?64�#&��ɒ6p��)P.\XI�z9=#��G�M���M��b��
{��\�ឝ�
SqRX����z�����veN#À��-%	[���h��O]�K����ׁ߲��x��P�*�Y�tc�ѩd8�(	G�_���~���� sq�3I���?�K�_�����K=ݡ�@�CP+�dǍҦ���fŹcC���<
�;�4c ��H��#Q���9m��٦��A_X�%�A2sa���kA.���So���`4\��4@d�.����܄R�1�h�*���ķh��7�a?�6�T��Y�N"��P7젚�����w�{X?	G��]��	��Xnv�b�2⮬7h*J�J�D���W���o��}�`������s1v��o-Ue�ͣ�|�,�﬘��*�{�A4eD�G�H��G��m���W��b����܃��i@��DimE��� � $�������M[rh�ﰒ���~�Fd	� PG���t�N�	[��p��b�7�x���Մ	�#�N���	���U����iV�U���H=�5�7�j��~vr��������ɧ�xܭ{��
�s1��>��+)�|Jg�C����,��VbM�/����ki(���&bp�P
������X�:�Ƽ����QYV	(2Ϟ���� �Ć#+�OE^�	�	�a���+�g%��r�4d�ƕh&���VQ���i�{��%XJ�e����|[OȪ����g����b���}b:6)T:	�=u�m$tvz\�U����B�T,FilyЧ�l���9�P����%;�ou���Pv� 5%���xW���s`7��+��2U���� ��>�PM���@m�ِ��G)����']���]���K;p�x�hF��u6�O�n%��0s�}�Z�ډIG�0�C��N�ۮ�A�׼�/jը��"�c�z"�>��n��l׻�J�|�>_�,�y�h̰ �	��z4|�(Rhh�v���M̼��H�� �Uo����-��i� 3��g����F0O�b�����'�a�T��y��0'N%���Y�X�Bv&Ea��AS�` �݇h8Fr�SWl4��d�9qusԩO`�jy��Z˸s�R)7ۂTDƃ�:���H���u��Le���8�? QdϺ��bHs�*��u��x�� �hW)s�!9�:����*���� �!�[����ỡ�$��.c]��F�W�H��A[ex����������qǷ$����E�?�zwN��J
��*"�5ι������S	��'a��2Y���L���c�P���Xߛ�	�!6��tf-16U~���V�����u��L"wEw��0�>���)��a�
x�pj��S�Ѵ����<$��X�R����� �s�7��|�M`��J�͛?���g��R~���Kʹ��HdX�����a�6�f;\��x���ΐ������W]�D��!@Ec�>�E����Ks�_��aQ�
�yi/⯵uí��q�콣�(&/��5�0���cR1��P𑕾�Z�:, ��xݘ1Ǉ���,a�25�F�$8
�??./���Xy�1���	��/SѨvA�����0l�HՎ=��Z����C����6呾�>�W�7��n\?`n�;������Ϻz_-R[~x���,�m���"4_<���%.A�_bE��9n�m. ����F��
��y����*��z�P���I���%���@=8�}�Lq����� w)�pU�i�W*;PA���p,������Ţ�Q�ߒ�y�lI��gߍ����Q�hZ��^T.k�M���2d�����%�ڷ��j���ޫEr����+������i�>��Ud�z-�n��5��y��{L��0q~��R��EB%s�>��=�B!,�x������I�yo����K�����+�r���-G�.(�sr���l ��"�ڬ���0��\�����o6�n�j���k��z���$6��:�Ͷ�L}_Ɛ�بY&��2}�@>Ƽ�Rb����o�Qq#�EY]�2����8+dq�P"4cS�۔D�H����ð����ꀝϧ�o)Qt ��?Ѡ�Sr��'M{'G+g��#]f2U�4����4��!p��(1� 8���ͫ��:\����Q�	k��D�q��{GM��B =+��19A^Se���MχN'�R<���V+����$�BS�L;;�PB�=�.b��[����C�ů5�s��5�3��`nq9�0c�V"���:��`�2�����y���M��t!g$⵽�$��?.�}����@������0��?�<Q��2�<���vg��]]?��-="BE�\�i���q֌�����)E:�c�`��Ó���?��$~M���^�lwB��_sW9����(�H��x�]b��Vvi%ώ��qi�%�1�ӹ���-/���|��ݽX @gTL�Q"�bT3d��O�T57�A��RH��l,ve�d�K�l��ߞ~�f�a���9���{è���m�ʳ���)7�:����O4��,��mųOy�9L��ە��e��"�ZH.2`���.�m�p4%�z����r�-�<[<���1���=٬e��64{-�0h�����[H�%��5���8|�Ȝ��-���Р���@�����ą�%�<_�PR������F��Z:�����f�{�iJj��n􀜃��{�n�uja��i(y[�]1^eR�΋�觻Ɂ�|~��r~FzJ�JhT��=����K�y����i����� h%fy�5��R�]�ܿ6i�bU���e�*~.������X���T�_��%�>wa���^8�F��T)7I�Fll�>�0�rwj)�P��Vk��Nz�	<���Q��I��٘b�L<��B�ȳ�F��Jci/o`�ȅ4��:A���oDH��NX�n{�B�1&���D��J�=�~�&,�:vB���D��r��G���E��l�����ٖ���ʯ!�gD�Ә�q�`�#o�:xj�0��N?�������G���_(�Ԧ8+�����h�rM�-��f�=��ZN���}�<jUk�:9_O��:��݇�����k��(������"쇔�M��OE�oٞ0!�vU.U��Y���$�$�K��hD	���1c�XCtsȐY2묆�����+�S9��^�ǶU#�_aW�:��s �@��>��߆97�Ȟ�f��r]$�8��8z��-�}\���Ƣ"ï]I�`dt�+�p��=��ᐙߒb�o�آy��M���o��!�+wG�ֲ����_ԯt�2�[��F�+�u��l,�k}��zN��	e��g��R��oG�3 ��[�X��ߡ>�����2Ơ��y�d��,� ��q��Y�$��`tR֕��A�K�,zbG��ݶN,��3�k�]R4�������Ep�W�2K��&2�[\n��k8F�,ccc�c�w}�n9Å5uuZZ���HP.r*��?S20h��9�W:�ɾ�����������'m�۰�Rɣb=�µu���	q��.�F� �]��D��%�;�'�T>˅�GM�;,�-m
�k�0��&�B��:���x�R�5�Kf��|^u��]���k���[��á���/���({.��m�_9�2���E���5~G}�'VB@��Y[�u�1=u�葵�դ=�Z�ސ�q�H� ҃�BR���x!��d�x_{�M���3�q� �3��������1b���W3+�� s?dMt�~yZ;�y���*��ž�o, ̮Ӡ]Wv�<�l�P�,�f����g����`ۀ-����<gM�O�E�GӚ�y�M9&s,S�jڤtf�H�S�;/K�g����YGw Ńzy��� ��S����RH��'^�c�v�kQ�t1A�l�
�,DaV�c�y/l��j?+�J"i�Q�2����T�W�h<1���;1���Wyu7�c�$�4���2�ǀ�����c�ʶ����'����̿����q5����_J�$p�}<����.̛;U�����p�i�g&��6>u�4����"x��@O:���a�����΍�t۽����7{�\�b7��X���.�����;��}�|�J�
�i����]#�|T��޲�����/�I��� ��쉣t0�W��ɏaE�	����H���V̟���I��N��H��["�Ӣ��A&�98�7�����%nE�FG�IR5x5-��
��#�[k)���D��n_�Qx�=��8(�+��n�zM�Z��=Jz
���v����-��d�����/ �;b���pS|:�&����N���tYcd㘽��Dd�A����VJ�rR�BW5�G+1�<�����T4?��͗\� �{�?)op4 ��W���Y���o"�q�U��l����� �;8p�=')�μ.�� bp+O��`�EO�Kd��@�jz���!L ��(� ���$��-rԿ�'�O��� ��-��e�k,]�0�!�=���*����[B���Q�p���t��Ė�z� .��L�,���tF����..k��;1�hO ��Hy��6�)=Ѳ���d��\)l������7D������p��kó$D�O��w�x�Nu-5��V�4�h�{�MU�&��M�H}��P� � �iʺ�̤����b�@��RE�������ˮ;!���n��	_�*��6�����m_���w��c�v�D����q�^���9�^���$�c������eɠ���i@a���.�ݟf ���5>�5�<Sr�.Ȫ��0O��Ok�=� ��F�e~b{7jmn+.NG�XZ��r�*Lz.(;�����v�.q>�o��- �<4�@��,|0�he�<�`7���r��0�����q�{IN+k�u��i�O�8�����V�7;wT�q�A��̙��� �kʖ�/AIEB�+9Yd���߼D������9_o=��&Z%#��e,|��.��l�M	�I�&Ȭ��g�L%�TFr��"BK���L�"�z�!��%	�
���ߡ�]R/�з7�C��dM���\L�쾐t�!�?Rj �9�r-���"��8�Yf�i>���ѵJ�F��Z݅�0F��w��׬Һ��	ѯZ��e6֚���r�dk}Bl���:�!�y���ճl.�Ε�̛��m��6��ζ�<5bW�FO_��W���ѥb�@��^ZF�Wy��!:������� >bV�xY��d�	۞
��;8�9�3!��H���<m"�чu��L��#�X�	P�1j>C3BC�[zF���p����r��(26�I�� �%Zӓ\B�]@�1��j���8OF������p� F��B�\$޼N�roɮ���\�_���C�r��&BNFQW���O(S!-�lv6�:&_^U�`n�ޓcO9�o�^F�vѠ/ @!I^f��Gc��dڕ� ���>����EQ[2T=՗�'�3K2�>Ah�<�0���5�%1��1^9�ҷ���Ǿ�I	Z�,��aX�7�!I�)RF԰��r���h_���dsoV�!~u��7g5M B�NZ�����"�M��-��5�q�t�iCO�*��Q�E���;H�w���|'�FJ��M�Z���<1~��9��%qӾ��cC3��J��2��`<�A0�U��G����
��֤��AI�HZ˲lJ[L# !���#���&YU|m���H�\��$�����"7�giU�&���ͦ\�Q;�5J?�uX�kZ�jb���eQ�)�Kc߆���R�獻Ǉ�p�X�r_˼�biz5犛��O��	)8�3% X�������M߯K��(�9�J�$�"�g枮Sa��k�8��.w��E[�r=��J=a��Ɨ��y� w9p�K4�2D?*.ubq��]�	g!�.���bd���2Ӷ�eS�~������Y�n�x�w{fs���L���WtBz�~�_U��!�1,r)�e#ˎ&�͋n���X0�(��O��X��(,a�����%A"h�!q�PͷO��X��Nv��_�Yv��&*W=4�W��h�c�c���	������՘0����CѝF��R^�c��,ѿ���"5����^�-i�u��"ei��6.z�f)jÃ4�/��s�lNw�c����,bzy47����箍Mv[�5�a��d�N,��M@���^��b+[E�_����U��F�p;�`� k�\!�c����u��Kqbv�B �_�uO�Q>��;�$~T�6$R�����C@1[im%��Q���*�m���Hd�0��>7[��ߦ�����#�đJ�3I��sռ� �|�kq_�&">W�&�ͼhz���}�m/�沪!�� �!F��#rc��%AbD��R�d��&]-���q�m[$���˧�3w�CLN���g��  9mt%��b���?�р����{�R�/��ٕ�/A�ԓp���D�����D�BCo�}���=��tԓ� i�M�
j�D�?6�{RM����FE���ʾ&0�l�[{~N���E/_�)S�7ľ��
�Ltǧ6H�q� \�0�:��M�^��ᇥaR6��?c��
D(,�G'ZW�'x�:jY��������Yu�3�ߡ�n�\:�r��,��l��sc��,엿��0���IYׄ�Sz�� +�8�����S�|��0�T'��B�B�ĤLq��hMeZK����G�Dk]Hj�TcC�#-���i3�*�C�5��� ՃlT�F�$����ܭ���7��[.$��nc��tɃ@R,�*�<�[0=99�	R�l��X��.`�	��&�Ӑ�����)+��w���`��D�o��xi�py+d��|��)i$�����q'�������t�k:eۅ�14������5z&����%�!V%����fE:cl���b��,��u)T�yψ��K��b�QB�����C�L�V�kH����nK��g]�����U���F���2�T6�ʅ,jY�b�"�Lǹ+.�*�M��4ϼ������b����2<*g�v�א �����%��#�Qf<��g#�\�Z��dA�2���+�f�1�>n�Չ��y�$sz�D����:�B`4�C o�w1V��ʏ>�$e�J-�0��?RSL���V_)���X'���-ǣ`�� "O�~QQ��|���8��DK4彅�` 
ݡ��P7�r?��=6T��W���9�ZK�ߍ�p<+���Ղ3p�:��-�6�P.	y��7lx��d�e�����j�����jw����ߢ�!�qB��?��<�}�c�V��V�̀��&�e(�1o/�Ƙ��#��4DP�S�G:�C� ��8�@�����[��cϒ�HD	�uUD�kF���D�#d��JA���p���?��@���l������4Mx��a�]o�d��;P�*�<�uf�U����`�3A+eS;BT}�Uʅo��mݤ���('tҎܥ��R�'��#�h�����:'����{�Ǡ�v|����ť�_"@Z" |�l�����R�e#��?	πEA+L��[���e_H^�k(�̕�]a�_\/b0��-n̚h%%��N �|$�#t?�<�7�a��D��_�]�.<t�4H
�4�t	H%��C��
)%��Р��tww��9����?��Zk_���f���C�Ҍ\��z�M=R��߱p����D)�<�s8v���S^��ql�8I. @N�B$�����^��Z/*�*.8�~�A�'�#�R���?#�l*�p���c�/��*Ƿ�@qz��I����7��ŀ��Լ���p��������o�˘���/�t̏j��sha`�.Ă���ER�U׵R\�@࿄���^��9����^���V���%�"���v��bs�/���E��z9�C�A�`v(kG�=��m��2��d��׊��D��	d�	��?�<p��0p[��E2M� �'�׭.V!�)���bad@#�C��N��dv��(�2X,��S0�\�V���	��ï���2v��b�>��.gR�uNy�'ǆ��Zt�BQ��7�}튴}����Ӑp����4==������b�"��N����J�+�D����fn����kFլ�"ל&;�R"���:��W�6�~�/��k)*���sן.���$�������T+'�s8� ��n_�%	�}®d�8�ٲ4\>�N��iC�#�Mٹ�@���̨�f*7��'�<U��MĠ��n#�ۜ?ޔ�Z����&�޲q��тVmԂ�p�-��)x�lG��]�T�h]�Y�*2���%a��h��fEw��h5�Xڽ�2��؅Ca%#��8N���d��:
�&Pm��H�\���2���a��"�y,D@_��gb�͞�3��bZϖb�&�������H����?�/��׊H��tXQo�Iu'���X�"s������|�#�}~�"�FG{c�"nIb�Y�g>UCy
T&���_��)�GХ'��[�7;�fI��	,��Y�|����iί�D�k0�۫��i���߃vr%t�e~�t5?t�x��`r�˸�_�\3A֛{�A8���Z��eͪ�����8Е�gz��61���
!���$��`Gh�Q��!�@Z��e����~��L�W��֌�s�<�z=O򸈐wtuG� mv�Ą�n��/��� <�W'3��U���Ȥ������f:�iK�����/�om��C���*� ��7Ym�֬�j��7�z�?�ug7>�6>?j.��k}U<�O��$����@��w�6�B ��[�ں������X\�:�L�@N7AN]<��wG]��9�hV� ��!���I��
�R���B�&/�t��G+����
%7����܀��Ѻ���z�������FD�eD��.V��=�^X� NBS�N���\�yo�N�*��U�������|�����+k �)���u^��2�)��f��#|=�PV�yη�C�>�l NN�@�x��0w�C7�4f@����-(�SQ9i$$ovNF�z��!���@�O�V��
�T��l�"�o �W�b����i`TxĨb�=��s� ���H�K}�1�j/��0�8�=ɢ�M����B���1}v�1�{��U-2ExEO��`�k+F���ȣ��7%X�Aw4����A>�X!�aZ�#�R�Ҍm �,K��h��)]%��
�E���k����>�d�7��|��e�����k�u"���`����l��c�IV!�}.q��˴�n��ꑩ*��K��\KC4�(� k�%�.K|ڟ�a�P��EU\�1���M�r��G �#��{�(��X����H��[��eϺ3�h�7);�U��=�����+�[5*�qtE�<
��S��ZJb�� R�[C�!�Σu��1)d*�hT���bC���'.^c���>����[U�ê�!��Ū��8����D<9���ꊺ,bV*\�m R"�m2.��X������#zQZ��y��y.�y����k ������Ië�ޢsRZ-�鸂ҧ������Z����}O/}Wzf�F�_�$/\�� TsW�I �����<����U���M�˪-2�T"2"}�3Q����Y���gG�U.�L)�9V~<��c��F`�������.�����n^��H9�2�5����R��q�	�S�����bT�'ƕ(�μa{V@�}s�?�k1P������F��U�����tZ�xSOM
!�aA�gE��n�UB9c��9`o��ޤu@��cY���/��w�OMhn�C}�L����?�b�
 "ҡl��{>�B=�D!J�a)�b�v�O/�f��Y)���'C�.g����D{t:�qppj��B�7R�h+<CX�����Eb|/.��r*,���\$ ��➫�0竓6���\�C=rs4���n�̔4~��^{P;��~{cݮ�Ɨl��3.I�*�A�<M�Psp���=]�_g{�ڳ7��T��fs/K|�k0^�	���&�ơ�U��	n�RQf�2��vR�%�%�]�\o
q���l����ʓ���mbO�WO�1Y����{&d�I��>���!@#v*9�;���Ak�^�\˱R�~$ Wrǧ���|)�h�z����14�mٕo4e�g���M�=�A�o=�Tt����zq�I��ˋ�4��x[�W�/a�((ւ��|��-Ɋ�,���s؜C�cTt��/ƺ	C��KiaXN�.5h�hQ^�{N;��i��v*��dc��I��C͛�Jd�sş%����"ᣙ���N�Z�?����Ϊ���x�	����/=�-�
����{�`!f��BWh���/SJ����q��#P'��$�w��l�bj�J�8D)��`7RRqt/�(=�?�6�b,[H��;��߮7��$ڼkV�Z���5HN� �u<��C�V��/���{f�H��8�h�s��ȇZBpm^��9IS&AL]�&V�0qQ�h /؛3#�@E�v��2�9z��8�;�l���)x��`�K��$��;$�3�yH+�� .ީ�T��Q\���� (]��8BB�C$*���,;��*��)A�"�=���:(�@L�ʹ��b���a[�J���u>��t�/�����j�YU�z��O��H������e'8�)s���=�,�.�S�aREY9,��aE=ؙ&�@��Ԇ�}~i_jK�9Fx�gm����i��D��k.4�ʛ�Y��w73�*t�+���'@.:a
c��kᕃG�w�;j����-&��%����q�w�H��K��2z��j�lޭic��G=A���&��(�|��6�(�}n7_��n ��4>�.�GCy�c,�L�Ӊ<�iG�l�	y�|y� ]��j~��E�c���!,s?��_O$
<�~��ڀ���*v����T�;�E�&Q�@�hw�����s���_��<h�  KΆ��?N�$Bӑ)fF�X��F�0�B�U��/���=�h����	&9���w��p2%߷�E
��Y01B��j�L�Ͻ�ԑl�c��t��C���s��x�w�����t"�-��k��x��Vy?��c~�}^�׳w@�����+r���&�z7�͗RS��|�0�6���,�m����k8�ջ[��z>zFN��)�4w|�8T�q��-���^�~���.��AbT�}︘�Su��_j��xs8^������d9�������q;��*�����@h��F2f�G��$MCL.��1�?hɟ��k=XN?�<V��� =�Ā9|���G[*�Y�Q����gsRz����C$�B�����^.u(D�&a7��N�	���z3˪±�+��w6�����e��Q-��r:�������/�5�����0�h���]���\�jL/�W�Y̢��ʧ��j�ۦn����b�4u$��ȼD/d4$�π�i�>�mG���OM�D������J�tw�X!o����B���o,�E��;� \D��=4�Yw^��l]�v,��փT�BDD��x���X?)Ӫr���}���� B�O�I��4�S���3���5B�J#Y'g$Sȏ��2� �w�د�c��c���0�p���<����vF�?m�Ȗ�\ʘ� ��s�|-䙽	)�s%� :|�y4�����49a�^E�T@y�:[�u��$���@�(U�Y�)�~ʷ-�9WP�o�%��8�� ���o~Q�7��"�����9�s��"��<{�[��1���(���M�� 0�*�k�ϛ����ub$9��B����l���
D_��*���I'��/�Q���e>h�\��ډl|�G�-��q��O�˸j� ��f�ve
-����Y�M���Jo9Ʊe#$\����y�D���0���Ű6�h��3 �S��S��Ř@�)n[�X�*<A����9m^�#~ުpv������h�B'r�O��K�a}Ia��h���ZU8C6[2�|��3շ b��:��gB��w��dJ@�����)��w�E���a���X���+��l��~w��i,^�F��0E4zy�����m͌���&���P�͡�3SZ��&N���{�ZÁ�(~O�mM����W������8ػ�D#a�9÷����e8���&f�dK� ��:�K3��
M�Wc���tI��	�P@ �j�QaH��^b��QZ̾�/��	T
�.]$���OaQ �z��l�$ mE;>H-�J��ᎧMc�o�����Ml��OǙ���7a[����Ķ�Gn�X���_ܙ�� ��b�.����UQM� d rY�����J]�&
~W]e����}���t{��7N����6��� _\����ҏ"=/�8m$iǵy��Þ����d�G��ɉ��@�d�� �,^��ynD�Z�b{}���.��S�L��N�ݸ�0�s�ܐQ�L5�%
��Ƒ��A�a�B����a�'���{,o/ݘW����PK���`�C�s��;$K�<�M�7%���Ν|4��Jd���}GnS֜Y�s1�@aC��T�:�:�"��r�!�⏵�Q�J��wʅ����@�R�g����Q	�����LV�R���믔����/)������~�Cg#�C����2b@ģ�@�P�K�A��&{"\��Į]�f�W�Q!�0Ӿ<2{�?N<�.� �0Lc��m6��/*�6��ע�?B ��9�A������&AJ��lez弿NG^�e��,�H������-�)�Ki�B(>,�e�h��y�+��e�̑�2��q�
�b�
�+e�%���u�f g���&�:o2u �B�-���{\��%Dv���NҨ��xh��t;��at�w�;ƎR ��z�O�#Ň�%�@N�N����au��w��b�"��C&����G!�h�^�E���Z7��`��<9�����秀�=j�o�B	=W֖[���Sh���?���3dά�X�����kvԗ?��j
J��CB�`��--X-����خ�V�Y�NP�1��z�oBS��H�7} t�D�L��.N�$H���өEP�i��Z�3�lCU<���)Ih�;Ev�,3m+�(Ԧ<Mc/�d�D'' J4�����T���Uj`��*ɷ�i ȏ���|�_,�}
��v�����1jP����\��?�X{�jU*�9�'�He~�4V.5�����m��*�.�fy���j-�� OQ��&�9�ɑ�N�1p�ʺ���8�9����$����.���Z�k��;�����GvY�cq���$����I2�>E��|h�3Q��D�`Jx���ک0�����ťfA�X��Ь��@�#!���M�B��Ǩ8��M�^�uOZv?�e�u̮�kU��~ua�_�UP�7��s02�-Z���Y�i��B���2���(��>�%GA�d<sJ�:��˷�H�'pݞX�����I�Aקc���F��*�K�����4��v��".֓ 6���+)�����:�j	�T45�w9OL7��=u�(|��XX�Ź =S!D�sz��2rC�{�dGYJ�?.�~]�s���=��ν�Ǧ���L�@��Ӧ᪰���DȔy����!:�Ui��@}�~i|6n�~��ݡ��Bq����9W6 �f<����I4C�c��E�q4_/Oq&��SO�~W3kǢ��S�D��,E��\����\Y��K{E�٨�Y������iE�@E��K佈���nx����bř�O7�Bl\���D�#���J$ڌ�,X����'��9��6�&!eNQ��z�����@
I�q�F*i%��9�����5���_�sJ޹Q�I�V~�c}�K#��|�i�Z	����3Ɉ{Y���_6s�-�[��zm"t�B�F#��������eD�".����_����`��M`���_8��7�'�s�p�_r��COK�:iF��p�^{�GiЄ���k�/�~ٚLP����YY�J�:ue؞���Rz3��|��6۰��K�Vn��x�(��;4<�Z�Vp�"���W-��N�/p��s!suK�#���՞�3�F4�Ÿ��8�r�uƉ���Ͽ�7����1qW�3�ݥ�q���~�M#�~�k��ʿ�ԫ��9Q�c;�ކ�����23 ��S�G��ܴ�9�;4WH#5��Ft9�s9< 0t�ظ��,X�]�
K��oA�������\]sG�:��V�E�q�4�-|����}6�bl۫�2����AOKR~/����Ɣ�b��U0� $|�/�X����x^=���$�CAVCN�A�H���\"@�-T���cz�M���A_ӥ�*搋V�Q�}x,��M��NF��vZ;&��1����˳}l�����n�A�M9�U�  k<!��<3:2%����pe�k���R���d��0М��69�VbNdR�����-���z\��|h��������iw�9_-rЛ�)�����}�R���3"FA��Q�2��7y�.�����@���I/WF�Ulu]ۊp|P�P�A�WB�մ �%֫04	�[]04��d��jd���"��>��w��B�����8���<�r��6���l�69�����Ik���CS������w~�{�S�m�:(�Z(��������a&wG���풂Fc7�R���V���B�N+�9��w5u]j�����La6,�h�G���&�2Ws�̍�b���a��%�F���L$k(��]�΅��u��L�.��:#�YJ�]d��L+�B5�� ӎ��y�IRK$f��x���_a��/%�`o�: �e�YQ��3����ϱm���q�h�)u���X+z��g�CJ�ر���P���_u�(����H�s{�4)�\^�=�ls�6���Ί���ݎ��.�z�L�+U���Z9���Y�1��)0�(d1����L�i.���4�����D��A�$1�	�������݉�e�v��>��C��
� �1�C��m'Hgm��+�;"",�0W���+���8�+i����qp.֞��`�wO��<���Ȁ��C�x@r�h{�ҔDтv�-h�Y�L�.�y`��i���I��q ���O�ވȞ�õy0��R_�y�Ju�<�k���)��u�d��6jD���/
���2�{>�5�_�T��J�R�]�w^��(��4tJ0�����ۙ@{ ������7�k�C�������~���s�d�
z�����X�-ƣzv�X���͏8dj��-VJ�i�Z���f����>+t�GDՇO3OI��ފ�I��5���	���߮V�����f�+�y�U�o�1! �#<*V(��j�{d:���N�K2�^.ic@y���-T���I�Δ~�،�#�M~�"Ui���n�{��[L'�����8��������!Ӟk{n���Jٕ�t͋��f�_S3�;p��m�R�>��E<К|5/#� '��+�������/���	�!uV!ߐ�4�B(��4�ͽ.2���\�M�䊩��t~���shL�L���m�ۮ7w����4K��B��;��&�f�s�9/���I"q�{�F��.�Y�RN?���o�ڈ��xb(�zO�z֥�����W1�P��hr�`h�UbKi�~�:`��\�ô�T�g�ɵ��Am�V��t��s�n{��t	INr5���;�%c�s
8k��#
.뽡����������D��5y�Y��@3�5��Ba^0;{�"��	kǵ^�.��[zA+J_j~i��ieݙ�v���X<�W�~I��'��X���L�[E�m�� �z�A�y����p_��GB�It���?��w�6ǋkY*4���:G Sm��M��uv�wψ��f)W��01U��K�������*��4S��>v@!�\��F��������Y������MTSGX�^R�fkK+vJ�r�4�_*���U����҉}p�)�K�B'��q7����bc�fٷ3Яk�@WI�>Se�/!�OT��.D:��Y
A��i0��X����1D��	�?tDR�u<��h�)[ȭ��e~+��T����)�xӏox���=�cpzsoǭII�3�/=0�����Gh}j����)�^��l�T��E.B���A��Z}��Bj��w�j��4J�i��<#]z�g
I��R�"��&;쪭����(���^���4�_���tȩ�<��F�m�ӕ�L�<�z'Q�R�\KD!JK�->�;�23�e���eLp��,��2�;{�X�d��QW���S�}ίi�T�o��7�P�'��z+c\�����y>~�r�\�T�Y^x��0k)͹vG��wӂ�O��|�"�%R!0f�jx:�s�Cױ��gwB����[K�~Ry�R!Bnh�С�����
(:O ��7�4d�(�
2�l����֜~��gyO�V�jٯ�6�j-��<%�����\6���<�`��'>��x�)�����	���V'!�R�S���N���aٯ�o�<�b�\�g�ƹ�S�"�����g��j6eSJ�����q�_�_���Q��"0}1�N��HѸ��Uĵx�߱��;9e���35�2Hxf"�UV�:���g�,T�lJt�Q�.E���}�j���m��r�^?tl}��NY�8�+�ߓMۥ!�W���4<UH��(lj��j�xf+\9�$]��+ò6��t�3�	��՝M���I�L����L���dB�k:k���q��[���o{�⢎��'D|V��Yg�t=&��|g��{ ��n$J�jL�K��TӼK�` �,�*%&;�K<p,�|�L��9b���uN1%����k�v*� x���P�<��;���O���.o$����vBr�z�3�	?�U�~�U��3k�U���!͸�\���|ucdf��ڭ�Ba�?�m!����y�c
iN�F�w|ٚ7������k��x�1�op��\/��k�^X]9TW+JUvL��T�J���6h���4� �U������b�mTT �Y�=�D��d^Gg�3#��qp�7��j��v�B����cT�+���,I-��с�C\��޷]Lh�T�\g������g�F�w1������;�c�(8���<c�{F%dR!?~�Li���̟�`�,z��l����U�˸��"$�k�;�����(O��꠴��P��Z^�v*�.�ܵ^����
��� ��dDI�̭]و��t�3�b��!���Vii|�*�Q��n��+Bϴ���?<���yGf���{��6���e	��?�B`�%��Iϻv�ͯ��������}��q�|Ε�M���}�X�P�F&�3p��l`i/���bI_�M�ջ[V���a��pNm�|�R֑
�wl��UU�c�
S�2U\~�{��N��^�n�#�)k���@ke��/��U�s�7��jb���;˿K:��,���v��_W5��|��ӿ�̏�E����(����к�N�'��p6զ)�
�_{�Y����m��$%��i�z#��r�]?4�]*i�)=�搚�	�4H�Z������q���7���M?_r�;���P���Mkm���<u"�Xƭ�T��1��e�y7x�c�(��ki\Y��'&��)2��
��e���W<=�h���s1Zq?��Z�<A����c!�T�ʀ��s-��y���]�4"�KQ�Ģ�(41jev.��CI�B	^4D�:o�IX��t�T�#������}V��o��=���!- 'y�>9?�ɶx�\Ͽy����cj��[Mc[��w��? ���^�윫�R:xx:���̽���e����l�(q�uj��"�ԋ8��^Q�/;��#;a�l*�G����Q�Fos��O����O�k�R(��Vmm�E����H(���dOi�} w����ũ�r��h���_Mo2!�<������<�J��S�K|s%�L�%��\�e*7�[:ƁB��� �t��G)��.�O�E4�^[�j��qf�8��p�Q(����"�z���(�/�뿿�`���_ǧ{�o�?��֑���o;�f�S���H�U�s$!��{jH��O�=���Q��Б̢J&�*ln*���mV�|2Z�e��ێ���ƆB��R�
� K�H�x�8T�QO�3��/&A���Aw�@��n�u�RD�\۫�@'N��@��-���(��c\S�8(���Wc?�l���J�b���p&иm�.a�M�(��Xbfr�)�)V :�d&p�k}ZX�z-�e;�!�/�U� ��̩�P�a��l;�㞙W�c�s���;o8oN���MI����e�՗��(��'�粏�j�X�6B+�Ǟ3k|g�D��z�'�+Zk��Xj���ۦ8���k{}��o��[jll�#Sh�1��C�@� �#ڂ`���@�|�~#�9D��>P�֮�,��k7�<_�[4K���q��"# ��"���8O��(�1��3]�8���r;|��SgSYT9��)b���E�pA�,�Ƴmę����Hx����M㵂�0N[	?���Ʌ��SEM齶H�9�����a�_��d�ø���<;
 �(QHp2I���'mm��F��!Z=?_)��B����:"�#:&�\�}(�
K�K�̳�N�!-�wT�]�,(Y�|�/L;�������ց߿{����&�������?�*��9sR{�Dt��O�f ?�5K�>��@X~����;&��A�lbx͗�%��R��]a?�����/�3��J&f�l����9ߝH��đ���g� ���!KLM��6s��)��G���F������>����} ���\?�z=����uQ�6�n��=�st9zZ�x:�4Gk�:�n�!!t�R��FW� ��vӪ"����OPs��
u��T���H�	�V��p��Tq@�� ����Ѥ��9;�w&�֪F�诙:d
��5������m,5��G{�!ȸ�c��]��_Š�?'6�c� �7�E�������1�lc?+Ʋ.Z*u��������Y��\f�9�?y�\�U;��>$�٧��2�2��h�zmpɷ_YI<pC@D��ʋ]���i=��/��V�����7��k��nb�"h	0(��n�)j畃�����L�t�J�<�>�?yǕG�U���"#f'b�ab+mw9dH��B9u��۹���_�����<��Ȕ<؅�h1`kݩ�P���Cj������_���qH�3�3s� YTᣬ-W�-mx���qY��6����a�.T��2\��Р,-��w-Y��/��b�{��Fb"�bط�'�En�z��W>F-��'{�cwsW��?�3
��.8��⢋��Fg~�eM��<��XȤ�=ʻ@���6E~�t����� ��t4p�*2�ҭ��Kƿ���&�m�f�C*���pH�"�����L���+K��h(��0��c�U���Е	@�dXv������͇��||�m�!�K���qgz�i}a�z]�A�����PC����W�c൯�F�����*#������k�^�?M�O�Q�������l��0˓�n��`#:1l`������Tx���t3��:�F�%��{ls����꫁�_���A���.^��2i+�G����ZKS���^
@I9�\�"��Z�VȬ:.�X�e+��JoG�;�u��9�O���ޖ����XA�x�@A�꤁@	c�/�г}�P[�/pt��Z�ښ��Tddd�]�	;���(M��0�U.QV�g�L�.��m��*Bw����,���v�&��ؕP�8I�/��i�'{����Å��ܽZk-c��\���m�B~C�*N���缊����< ���5r��O/Uq,Dd��+�o@�/`p��+,�qcE��m�G��JY� P�F�o�j��][�o#c�af&�u�z�*�^x��JO�6���c� 1:`Õ�{��%����b��6���!��{D�Q���aKOs��� ��ڙ9Q� *�_U�1d��}f��p6�x���S�D`V��|_�)��4�GޱIh��9�x�6�^o���ow�_RY5�4��}H<n�������M�$�~����F�����>��Qپ�yÔ���4�ϋ������Lv�T%
<�8kP��iX��qFsyE�Xd��%�� ���/��V|��<�jado���)G�ǌ��,����5]�ؐ������xZ$�A�Q����Dܳ76O���st��gF@�-�����z�7Y�Z�֒~���n�TWg���;+�C����ŋ^)�2����ɬM@	�=C�B��̢����}ô@=ʆ*>U�\�ٗk��7�h�~0�N<T�J�r�����\B8`ni$ՆD����ܴy��Bz��@���J�Xf��*�r�H�����NJH|(�}�)a"�<Jo�m<��Ze6U��uCM�h�L�U���:���:I�A`3�;v:�=���0"��ػSՑ[rx���*"W��'��OɌh�e�!��W���U�:j�=l���DJ�~�m�B����4���p�BDM*��f>���:u(�^v��#��s;�Ab�������?KOKBv����OS�s���3�u�ėc�r���G����}^~^��+b�i+�	��?��9uo���e���4YW!�7�j6���s�R�>>E��Gl�f���ZA�k��y�d���q���A�Y�KOg@�	����K�<Rw��D�1��Ƨrr�i|%\��� �Hπ=�:�b;�ei�8H�y��>[��/���րp eϓIA� 5f��AĈ��7��෨� �؅��'����{l|��������=�0�t����ڶU���r{�����4d����4#Qw��W�f��ᖶ6J+GR�[��*M�)C�f|/.���u�RPp��:�v�lq:�'�F�n��}�a\�tE&p��P_o�m��q�Ŋ��C��z\m��R�e�a_��!1��H��0�ժ~3�*����I���f)�G�hX���0�>ڒ˷~�]}h�O�e@-�3��b|��{�t�4���4���كo�D߮����d�ɠP�G2���淎pמ����)}��!�(?��L{!f'�"p>��~�+kf��z�(�Y&Jj3j<}r��lÌL2e�Z��gɬ��c�q'��)�<j)��QQ�x���n5����}�u���@X�W��G�/�Ol���^w�z^W_ԟ'�
غX�Ba�D9z�2֞_���������}��"2���Z��vI��d�ѓ)=6�M/���p>?�O�و��cd����Y���m�U�V.�^���WH�!�^2�^�=��*^�s��������〇��G*�fI	�_���H6< ]�P�^;hEn���L$����?!sBy4���ں7q
�7�c�$���4 <qj�[��j�MV�5W��i�wSӸF�XB#�2v1P֫�����r��Ɗ��;Vg�� g�ǳ���G�6�'�F֜��΄���®�11��� Bp�Wr�[�(�6-�4d�ꍀ`~Ը���59����.Q�}�H�L��1$���D����w&�BZ>�l����q:;a��AD��8?f�u�<h��^�B���k�ˆ���JT#}�Ϸ~��o)jj�u����1P�>��;!P���L!��D�۬e�Hn�T҆b-%���sE~8��`��Eh��$�:���n��\��w����Fۍ���
n���4CL�t��q��:߬<�=���x'�fA��\�+�*؝���z:3��â�<;�a�5�οa��;�S;nf"����g��_��!��5y���W5�Ψ� Y��X��
L0r�@��q��`���Q�NCh�D��x���}��W<���sS>M��,�>[U��Fng�}v�a�M�O�h�����Ih��tq�mf���*Bo�U�45���S�-(�z������:��-vM�������b{U'���m� ?��M�&g�'���;���r��Rug�`#,i���Tpu$�"���|�݈;|�	\���ܯ�����z봮�I�c�Ō ���:�?��S8(��U}���kxc��p�籬?K\��eN����l����WJ_d�pa�4й���b{��K-B2������O����1����?�>��8b�{�\'zu�ĹH{�����8�O�/2� =ҙ�~�TG� �(�L���:�t=�
/U�sW���a65}�v�ĭ�>䛚_�^���:�V��5��ʵޫ������IG}.��F����}�_n��ŧ�;�Ɖ?��Q!R��#$�5k)�WW����7L�na���N �񹱽��%3ق����� �B��ycGO3{�HӢv?5)����K�r��L$h9��)�Zz�<�_���*����z$6��ޜC�ć:�������*C���?���c~D*�Q'2։����8�'p��2�>��~��0��u���/ 3���u��n�5�S�gw�a�"+��X�\P���h�ɓ���Ծ�C�v����	Y���ַpxN�D�
��']U�j��S��/�niz�ğ�o���E2�K	aXф�o*�k'��￐�BԪ�
����M�斡�5��s�gwZ��%��U��E�<�ms`�G�R�x葚h����$�?%��pN�*X�#����]���F�dہ�QA��\l�aZ���^ϧ>x�B^�[o�w�2v��n;�:˨�:#G��;�PB��D$h���<韦\�-����8������m~wׄ��-&��g`{�n} ���n���4��q%����z᤻��{�WE��-`{d�Q�Ƭ�#*g��<^鱚�l�әl�u���w��~��snNǵ�2Y�GQ�ʃ"�"w�&Y�����7#�f�,84��'�bZet��W��"��j9� �)7�FF�r��	�����F��ﷆ\�7���B� (X��.�K3�H�k98�,��)���Ⱦj��B�-������:˷��HZ��Z�t����6���(�d���� ���N֖蟘0����������
v���:�D��3��8��f�_|�����r:Iv��(��g]�w�~���!�e�+EH��8˙H�@�M���j虄 �(�Pp1��O���1;�O���K���+F��M�����e�f�GC#�`�5�!��)�$�(��J*�)(���a�YY1�H�5��W�>T�/ �%p��^稐��2��<�u%iOC�wK!�
$��&�ωM=�nr�i^��Ie�&��S��$W�R.3��x�a֮����,Y���Ɔ�nM{:4�G����J���2�Z�k�$K�v�݋S��=He����Ա�^�Q�@���3C`�}H��8JF5����K���DKE}�O��j�_u�Q��|P��!�$��`z{V�I�W��������Ә^������\wl��8S:�d]7V��;_فl�n���|�?_/�>5m��!��p_Ya�T���2ւ��}.s���������.� �4��C܀���,���F�lql�ɱ��y0!$���r�9�yu7m{���v����vT~b(����N1o�7gΙ�^�Z��{b�$�5�v�Ş~�@�x���%%����n���9�-8���Ҳ�P� ��0�'����oDɻC�f�����=�-B�(�	��LT��Ή����n��aU9#׸�}�<8��-�m�=tny���z�H�V��+�e�'bl��Q��U�a�,c�y*o�.]e ��oÃ{ߞ�����H�0���U���vH��탟Ꞓ��D�E�Ոr�*T�t��Q��*���
��n���~e~��w\�����m#ٹx�=�� �OqOz"&� }�7�VN�9���?�)�ļ�{�\�@j��rR_yh�E�
��Ǌ}ן+����?Q�67x�VW����<uv��㩿�F�i�B���.b5��z����x�����!����a�.ɡ�S:%$��[i��:}}������3���'�Zg�/�<�	�J<R��̋Ҿ��;[3��mP��I
��k����e�5=.9l�[� %#?������1PL�j��/�v�a�N��8�.��1g��;`<���-�1:ݱۧ��0��t����?�e��7��K�O(I�h�l���A�~R�F��7��r��J��_&��G�,�*�;?�p'��k�U���"��� 0m4�i�I�(���h�r��6��U�Y����gxu���8���Wt2H�7) 4���48 |r��r�Y��H`�PSo@���Ē���� ��gxh�:!9��f�\�sn�7��ᇋ}z2����s�l��u(�!��Q!�K,a"�F w¹��-��*�z���l#7� #A��ϊi�(�ˡ'����w�Ԛ^��B3�y���Q�ٴ���2�,~�G0/���+�FJ��wҟjYЙ	j����E���)Y�X\N<�.�c��� Ԫ�E�G�N��2���1���}�1-�#������~��s��<"!�>yC�Ԯ��F
�ײ�Q���ߛ��{w�z~�g���(E��Β9�[>�����r ��_�mʿ2$H�~$�i%����#��Y��U
��Z��Pì�&+��,ۃT�]<C��x��,Z����J�ȕt\�P7'��%B�싎A�(�+�?q@A�˦	��>~rV9���n�!�?���[]Rp?���]��QC�	QD�0!~��0��s����k#�$��\�$���
{��Y�%��뛛/Z�Ӹ�"�B��ϊAh�j�蟶�8Qم��R�u��+�<zM}�Ff�,Cx������dx"#X��˃���s�p����>l�Z-����K�e���������LD`�(|��HU
�!Էhpල�K��!�&��4BRY�H.Ru��KwX@Y�������v����mD^|E�x����(<�<�������װ��_B�.S�q���+Ȗ�g�j$�@Ϯ=��8���}BB1h�=/�G�ߒ��-���y�@�٘^��|�u�F�.������G��-O0W�(���'"���_�1j�͏���d|&��/�1�����K�%��2c)����dO ��A�QP�� -��� T=�3%~at�4��B|�����E`��qԷ���\�t��l=|�II�T���(\G�@�RC�^}��>6s���&d(3mu9	�y�(��d�1���h���6���r6�W�腥׏2j����w����gYA��Ng({?V��H6mz�-���"�4}}�[Y�=�	��1����|S��rR��M=�t��b���8����)� ܎�`���
�g��]H�󤤄q�C+��n�2�
B��"�_����ю�69����
� x3`ЄY"
mMqo�x��"���Mb�H�+�E.���\����<0��a�m���l0��_�}I�"cM��"�+~'�A[@��o�!˙�*/(����ߋ�S� c����*�5�.��;���|�h��3��7æWҥ°Ň��yPz��3���Y�2*�4*8�Ϳ!�X��@B��v|�h�s ,UV�廩ا�� ބ3!r�r�����Ƙ+aC����_� X�������D�.����7��0��`kd L9$|j�"g��矁+FVZf�	��	p��C���3�}�� ���Q���k �gH�P��q�����ޠ7x���KqֱC�mCm�?'�(��+I���6;-�J�!��;����2����_r��3tl����� ��l�'�;Te�8WR���T�'���z�c%�1ަ �@P�X�Br�γuL���7�>��Y��(gDɤ6�cN�t�=��X��x����I6����Y|���	�/\��t37T���d�v7�����C�^Im "�������+�_܋��*Vg"�t�(��[��+dՄ��x&6�|~���Ӡa�.�LA�F�&�Ϟq��>M�+�?�
a{\|ьj��DI<�O?�{�b�#�9���v�+���WO�(�Lvn���������w��	d<��犸��*H�Kj��}A�,8	fG�[j�ʀ��?/l�ӑ$��8�?$�lsCpxԁ�Dx�u�?��EΞ}ҩv���w����7��Dy��9h=&����Μ�[\�!�-7⣊��t�@=�S\!d�|�z�q��%L�?d�G��!s�� ��V"�[�}4"E���d��.mʋl�p��g�i�=_�����BH�m��gES�-�ddU�溭�t���T���s �>�#����f>���{��.h��'^���*�C��N��)�	(U����y�18�+b��'�`��*�����F�Fv�n��~p^�B�M�Sc���o%��M�s�$Jvc3L�#2^�X�)%&X���,+�����X3H������ڡ߱��������a��S�>��(��	��@�u��Ih ���p(�#��a�}g���7�M��Y��[ )��Lԧ�s]�zĝC�F�G4���x&9�}H��g�7�"`}HM1!��ty��	�ߧ��~;�W���5W߿h�J`t�������V��M��G�<\�.��0�7^��1�x%�Q ��~���A�f��+��׫�G8��6�~&�P�6>�`��D��A6���iax���T_�7�d�W�NM��!�L�o�|���(����B�C��-S�P�RO sjA$�0C���2F:�����u��>o%VVW�4�/M!�i�V���g%���<��C�C�M�5n�Z��� a�=wo	6��æXƕ��A���K]��^��_YPՕ�E�B�;�'9: �#BX�gO�L��j��ׇ�^QE�WQ_}�"��o���cÓ�,߉O3@]��1�4���8�;��LGK��v|j��e&%h=��m��)���t@AjMR�՞�7V@_4B��s�����-�:B�a(O	��@E|�I��$EA!�^Ix�t�/�7���ڭ��H@YKQ¿���3�bx8ɦ��Kyy{(pn������4�Q��<$8����E��� aâ'���/�d+�$����@�	�^gko���7������q�x�(����BNK�T�rm
/\a��¥��Ym�MH���4İ ���k�H׾��8A�-�ko[y�Hh�(б�B����1��Hu� ����2²��$�:��GNH�»��dt�R�UB˘�t����Ϩ��h:+_3��99]8�P0�Pi��X�zs��g�J2�0I�@��,}�-�-��wRSI�T��5���V(&��ɘ��dh�-H� ���#��mJ�'	���H��\=.l���K��h�9�jm
\+����6g�/?��Z��73!��r!Q�����|�(�S"����ǡ�Py������! ���Oǌi���sK���B����O��a ر��X ܐ���`�|à���_p�û����Gϓ�)����HC�ad�����SW�ţ]�C$�%#�����ڔa��TS�k��Ͼr[-q,_�kRQO�xj��ۭ�B$�E�to�sĊ.�9��3j,B ;�oH���}�����!���z�`�J|o�!�s��e5�d�e"��	��#�L��0j������{MW�xםxK�	���=�P�WC4j4����*��qIN�pgH�t���j�����p��<^�<�/@�=�'�K�7?>���*}j�ON4{��TU��Pz�U���yu�Zݐ=H�u?-"d 4v��14K%��.����(���j���|��2������w�+쿽���͞�5
��ށ�-�?.}�;�ɵ�W�b���@?�r�����C��Џх:fT�B�c�s'%=K������ȷ�a���51�;\_xΈԤ��cw�d���k�WOt��YY�nI���.z�͠,�J�kfo�x}	?��_�0�`� �K1i�)_�� ��tɾc�椐��-��"��G�hNI��:94K<a�?hß>��
 h
�!bK�=��(�1�-)L�J=z&��>��4����^i��WpT���r醎�k�R��;�_��;�X� �Z	W�a�Fh;Zޤ�r)�M/[�@��������8\D�����_wQ4w�.��o ��9��=���u��au
]U߯�o2��#.)*r,p�;h��ayZ��[.��P3E���v$�/��d�}KٶZ<�A!߃3J?E�G�w�4y�XL�%��߱0�0[��?�v��D���w���jSa뉐ω���TsQ&��
.xG�I�ǉU!%%�h,{����Ri�C���ɫk��|�1ȵ^�O �δ _���,<���� �,eҺ�B�%z�y��y=[��e���:�M�!}Pxk�z����4=�G�޻#���5��v�))�`Ac[:j~���͎ �B}���s���	�p���	a�,�:���FeF;�F��2���4r�යi3����,5�|���8^�MAU(8�k��3P���vW@K&�u5��-MW�\G�H�I�\��D=xd� l���3�Mg�/|Z�Q��QǾ���Ќz"��$�R����v0^�og�Ш12r
A�_E���C�N��j�>�� �a�u2��9v�\#��k��!�ҙ���P��58&:@Dp�M�pBR~Nr�v5}�����U�CC�5��>+zx��
�8h�:3�xF��	)a�D$#
��ƞ$JKI{XP�[f�%|:�7���`��:���o�¹�M�p�Iګ��ɓ�g�j����o���-����g>%!ӈ�)��,��3�<JlS�<��h爟b�v�߰F#���NwVx�s��i%2�D�f����� x�߳	�m�05�H�-������7@f��J����#,��"�������7����8����H��F(*���8���PD��W��ڻ@��޽�Y�6�+�
lp��Sey�R�z�6@����$�Yɺz]t�=c�;1r���W"��Iۈ����3�5+�z)�Ĩ�gO���_		;�_�>�Pzk��]��~l�=� ^`�O���������UrZ,)��Q�_5�h���e{�������T���8�����/��"���.:b�.[zC ��J���L�֌�׾pn�2d�M��.swd��L�G�4�t%�zi��\���k����+3�dF U�M*�lQg�r>��_��k��)��W���4��ғY�}���\�g|&�ETqA�W�������W�܎͘T��f�Mo3���N\�"0"��=gY^[�'A�47@�|"dr<��}R� κx�s��k�p7t ���>C�_mn.��Ñu�٩M�e&�� +���daT��vF�81���/}���.��5�DԂ����� ����ch��21�����oKpU����%�0�s1�_�m�i	��"��bZK3j�%�{3N� b�%x7{ꀼ��2]�������t�S� W��\�^�Z�E� tH�;�*���0���F,����P�������ٽ_s�'y�I�7�Xh��$}�`O�1<���ʞq(�=O��,`�L�N�X�z���>Q�:t����D������cS��c��8T��׿�ʧ	���T���j$��L�	H���J<��³22��;��T��������Z�Є�1a���,�qԱ ���_oS�vi1�dV͋�8���Fr��*NtOV�q��-���((���ｅ�,ٖ;-]],
F���_m%��-痮�Q�X���<�m���t6���TɅ\e
�0띃�%H�%��Z�?4S'�<��E�ѽR��#$��+T��|��Ģ��@eS�]��U,�D�&�XN����,���텕7�9 �tB��.I*�����l6�ሳj2,��[�Ed w�$Ԩ���0��wA�^G���x��@>x�]��:�B�J3�QF��A�%W����pWo�	�mI��lwd�^��%F��ܿ����6�0H����C����ԑ@��󶭐�DQr��Pf~��_v;�Y'�K�5�6���3	&��Ewzk#hI��V*�#�ԩ_y�x�����ߡ�!vQ�ꧢG ������I)�%�K�?t�z��QI&��v�����FabIH�z
��Z:�Q��5�b/���-m��؇	u�0芄�7��8�����/"%�E�թT�G�#�W�>�>$UT�rP�
��cxM�}��[PpF?�|IwA� f�Z�+o�pz��)����ԫ4P��9�@����s�-���C�۞gzJ�ue�~#c>'%�=C�0@������i���6�А+�u��܈}���|#�U��&[SG@���a���
�xnS��I[`#��g"�4/HTW�'��^�R�����*�D֙��J��� ^A�C@mS,ǜ0�⇉������������v��"6/MpH)�� �ZĆ!�(�&$��ʑ|����ˈ�B[I���Ұ���F+�a1�߼�A ���G{o������ruC��E�nd�D��0��Qf�K鸅|�g���X�[��GY�����k�D�Ƿ��RG����-u�ј���=�k�H[�3�Y��R�
Z�������Y��Hؠ2�� ��[g�;��j
A�9��\C0��M~~+Y�ac�����_��7_g;��Ā`��`A�q�B����$Mg�WA�����ܔ���R�{MIz.�ٖ5�b�at��0����S*ɰU�0��Z��N|���@��'r�\NH���ȕh�oi��-�ʛ)q�OA������`���r�"'EEhZ���VqBk��ldm�Ѓ������,=��+�xT���m�w��7�`B���\�U1���2]�t|�
EuTƻ�򻁩�"]_��3��ªBX&v�A�=����z@��d��	6���,E|Q��F��%�U�:�x�e��i�6i;i)l�͛X`��.t�w�wl����g1���ϟ��x�W��N�ׁ4�)1��]m�}3wYM��5)���ސ�������@�<(�E��3�V�g�~,JK&�T�X�*��7��v��`a������Y����/-`q2L̓��a� }�%����7�aa8abbG�$�D�c>�JR98��5�;�V���"1�����*��7�C�e�=�+%
�,���s/#b������bY
H}SO3�$�����Y�X�իg�O�y�p�r4���y����4�x�|�=u��{l>ճ^��qB�n"/�A����ٜ��y�P��ѠCV��ꄐ�O�ލ?@���#��r��6]g��Ϧ�2����.��E߱�T������'8S���F��ك�P�y���G	��'�f��a�8�	�y�ێR����b���[:\2�71��6�­�vs�0�n.o�S�>頾�ϓ��m�|e�i�"Q.���v� a���n�>��������z��NF.��_����
j��N_��x�ÜW���:�d�:1B�!�#�o�u��K��G��<k$���b�+�6wB&�7�\C.-�ʯ8�Se�^&������U1T;�؍e4�����5[ �*`{ٹ�� y���
���RC�pK(��G�?�_z ����}�'%%Ea�@X0V�����i �n4�]+�3��$�����H�W��Fk��=*|2s��1��-8�r��0��ٔ��~L�*��48Uti���t���Χ�����jI,��D�xS}�{��[�O^K]������
C����6(l�Y�b��*��,!@�JRX��I1F��+)����q�+Ğ�h�����jM�R�";»,�Lra|��+�S���1q��3����u���j~������"�T�v�E8a: �Ȩ�$߼]��{�&�����rc����n��n`f:f�Ҍ��/?l��$�20�(�f�͸��(�����h�E�_(��(	꘺�%�5ۓ �o`�CzEi������j�5�2��`f���ܠV#M]p̟�s�)#��*ȵ,F�GޗQ�����*�0H�YDzj�[���ݼ ��I�h �R��EJB��O�E�}�1_�Bl���_"$?�Rļ���p�%)��ζ��K�~4=��͝�a��i�̏�t~[��'K7�68L���4�'S>R�o�x_�Y��6���Ap[s3|pUQ�=�K�`����o�|��~�s�$�P����m3�sFZ檻�	_����u��=X���|��x�o������������ye���m�x	��TZ:k5�Y�(�
�_⊐���|ʹ4�_-��&�'��z���f�����|ј�(�o�L�[�0�}��jYx����{���b���/9�.��"�	���u]�c}��ٌL(���3K�=��3�}�X�r�G�y�<p~�Z#.�
���4�D��L�^�&�����̬���M�h���3��P:[���2�U6����[6���uvDl4���?Y��Oj���@��袉�?��YY��T)�e�z�>�%UE�#��H�x�9�Lf� ������D��q� Q�!T�B*a s�+aDĘ���6}x?�+�q89��믋��P;�	� ��Q�t'������7{���n�`T�TUE:�	m:.'�i�^/S�[
uV��K��<7;ү`G�HYT��j�t����9�̺�S�N�M�}���P:qꛛ�l�� �B5j�������x9LY��ATƏ]Ls�sgk�����8�J,7�`��=��S&�5��$��	#�1+�2&�yB�6�B�z� �]��ىZ&�Q�9\�����"��Ầ��9HZ�n�m�P�v`yfׯ9��T�����e6�3'�u$F���>jg�/|�	���l��]��xfK�ݻ�Q_Ц������7�~���!A��v���x��-ə�E��D״v��y���3�E�Q���i�x+-��F��rAJ��B�-eb����T"��8��8�[D�Y�ZQ{�����qT��0�����2D����h�\P'����<�pJ���|���Ԋޑr2Y"۞�5˔��v�����$�S�Օ�N����.��ǥפEo㶛&��mB/��,�P	Ԯ}�Ȑ���K��N|\W����1뜤K��W���_m3wr�{���a�CB��;'��5�����p�_J ��c���aF��)�[q�e?A�ب<�����tn &f�t@ǓB�;��w�ɾ����3��_����ga�~�o�>*���q�M`7%���(�.s�H̅/y^7���N�1J#i��S��'���*H�9��I&ץ�خo�q�j_6u�p�}tZ��[H%�jsV�<5���g�MCAiK��|W=* �UR!��Y��­�����m��a]�7�����K%�w^7�b�)�EU{)� �������+�U,IB��<]��S�O�
'�<V��3�6��c�e�E��29�"�&ih�>����G8¯�~��-���OJ_!DC%�u��:����.�2�B�/�t@�G�q���gu׿';(�k�F��[�1J�P޾&�(�%�J��7D,惋���u��a��01��QB�Q��5<?��� ^�-fq���a�qy�j5�~�o��6W�6W��k8������k"[��s���|�;�?����oc���Uқ��.o����6��al���٤���l���F�uA4�Z�-gqۤOL�5�x��	�i*t}(tj�-����1� �&`�����Afs*���v�z�c�'2���
�������n*/��g�w�v�R�?Ч�k�j2^I����O{���Ō�mO&�U�ʵ�"���9���,ds��1������b��0���b��I��EΤ�=���i��i�E�ч���YPWn~����H��K�q�Q�	P��֚=�W-t���D�d)�҆��Ș���;]�`z �
6�
�[�v��{�Oc`�Q-���[�]o��j��q�v%q�4�tJ�J#]t���(��Z�������[�=m��HV����įjG6����W�k��5��e��m��Z�%��t������FP>���S���]��]62נ)Y��i��'�`�ŋݚp}�ѫ2I���nj��l�=7��ؐJ�~{J�~��x��og�@���v��Xk�-���}>_����u��l҇a�������� 5-��78�����t3����{h����΁�������a������$9�f~*"�8r�e���=[�����k5�;�a2��6��(�WL;�A���I��-%�{N$�R'|VŨ��������d�9����py%�P���H�e�A+�*:����m�~�?�Ul�4�en,����k���-@��ú��NV�t�%������������{�׈;�)⻧�	�y����pYA4'��&�(Zͧa��cW޼�f-�U���GC�����4�P�����u�8h��J�i��4\��'�j�����_Qگ8���=�m�I��]�G��r�ssd��S[ʋ���(t.�K����si��U��X�����9_�Zb����q%^@V4�b�s)�Y�0s�0]3xEK�G�^�^���F���X�ȫW݆�C�@^�	V��]��+��%Wou*q/���ו�6T�YO
'����G~��OKI����|i�&ٮ�N[=#X��n��^c���y"s

	�!��<H����c4�i�����_�l�Y����I���&����[|�����?���`����Ϻ� bF�(|����ͱ"k5Sl� o}�A U�N�V�R�g�z�n}C��e���1�����Ɵ<*'e�D<J���Z3Q���~�rDZ���S<����
.CaJ��o���5X䀐��͋�����ER�V=2�]�56��'���`Hg�"Ub�1R�èq��ə^��ɻ�ϼ���v�&c�I*`H��oj�]�~W��y��>Mv+;E�3�e?�/����i���&ñ�f���U\�_T����2�_���}��.Z&���j���_�;$��޶��J�v	&��`�ҲNƽ~�K�V�C�FYKወ"�`�G��l�����ܸ�.fk�'8�2��7p����i�)��%��W~$΍Q��a|�=Z�TQ�g�4������y��O���L�D���{,7-��y�9A���nZ(�$%=N�r����>�Z8l�}���#�&~^�/![%�+W�n�K;[��?��4B-��cx<J%���
��YdUS̳�펢�����I�a:��*>Z�;��$MԌm�Ñٵ!�Onw����?�A{�L�{�]�L ��>���74<PO� 0E�FL±S�@��&��!k`�3/;]PP�6�/��Q['�2�+/dUf��c؍)�M4�I�hN��#�0���~��.�������~lPSY���=�, ��5�kC��ᖯ���{ŎDg�΀\�~����R�7ŹkY�b��!w�����]�i��p��~s<�����5AR��Ay����Y�#�V�9���y�Β���=��Һ�c�m��3������¾�CڨEln/CA��C�o�H��k���</��?�pI��?}��6����e*����ݷ��_�q���ף�E#����o�Qx�5�l9t�n��k�^��gL
��^�!��e��H�����UƢq9��O�-M�j�7i�Vg��B�y�`%�o�u�������
�����y�[ʱ�̈`��}�)D@x���uOhuf���n"@��$�C/�A��RTd�3Y�V\O^��9����w�$F疨|i�-���՞!���a=��v����s�m]>9�6�҃	&�H6�3�ON��`T�$�_z���|�9�G�Ɩ��Fէ+ }��S�a���C�Yk̗߿
�CtP�'a�D�9�|_`�`Xl\f�A����jIQeݘ������s��N����o,�_Y'�q�����`����<�a�zΙ9�9���Hpg���xr�JV�L�^���qnל�jrc�X��K�=�&E���r^�i=�o�v��Ӝ-�U�N���I��ۙ�aHl���v�m1��W��*+��*�L������i^:볛�n��۱���5:=[��EM�Vo-ԡ��3)'޵=��Z��z�ú�}��=&�C�"�1!��` �+%��0�����R��96[+g~A_-!q�� i~�c�@�~~�Q�(-6i�'#�4��e	RW���ՙ�ǖK�M���o��������;}4��E��#Dro���η�p2�a�+�p��j�Qs���C�	�
.�,X�2;`TIU�R�XM�LA�����{��qS�Rm��l�nM�B�1��x�|���_c��j�<A�n	�>�w	���N���ds�^@*��6��𵈐��.LW�P3��ڶ]G�Ҭf�����.�#\)��.���t�K���i{=29;q�cn�/P�p�A��-T�O�P�����_���zE�H�45�8n�LETݦ�=-��ؠ���#c��L5�Z������4��`o*�qTgBe_V�*4��x�1'-��a��+l&������:y��pߜ����=��k5ɻ�햠΃�	L��~���>��i�U�|c�����������c��qSj]K���r���@~I�8c�3�2�Xd�Cw[�OF��R+8sp���J�%5y�9/�8��F����<fjF�&"��pN������m@ro
U!�����r�Y%o�}�Z��;����U㘙�K^�Y�Uo��׹{n�ե�J�|�9�h2��3��/G��������<[�G��<&\(r�4T����'��qR!J#=��)�F��V����ݟ�*�o�����h|W��ѱ�Q�D몪�û�#b�TTTv�����z���?*�\��m��ݞU1���i)�t�S�5Pե���7l?��@�YȚr�p;�[<o;�~,Q_�'�ظ@�e1�s�z�vەj�$�Z��S`�}�YW�@�\MR�X7���(ĢO�A��G�{Ng��"@���B�;��ʪ(`$o�Z_�(�jgp�p�V�μ���y���>��˾~IJ��d>������1*�y=���WA�T��i�L��Z}����9�񇎤E�,'	��YY��}�<�"�!���>�������xH`��i����9M�m���n~�9�1�w��m����ǯ�GUt�&ԛ�4�d3.W�c�o���b�X��F���Khj,�n䶇�YkU��g�\�����3O����	S���v����SS��a��Z����S�L��Ϯ�d���?u^_׵U�Ȁ�(�@�:A�����\Q����i���W����}-� ��睟�����B[�G(�>aQq�vُa�Xl�{�E2�3#�o�y dL�xK����p ��d�d;6�k:�dL��'�筃��/d7_7��;!�qUusv@V>��m+��	K[�,���a�"�� ��f�z��?��S�΢15�t�"ư�5���(�%A�I���5ߨp�"��S��ᬝ������)EܞXt��^�������/�n^E�Xx]sn��݁�߰�����a�r��)q��[����<�.�S����A���TqwޒCB[��>���|��d�&�h��Z_����(�c�5
ڍ�r�=�:����u��b�
>+˧���&+'9���
-�F�*p���N�˽m�˫��
�;��A�_���rpnbOuc���˧�Ewm'�1�rGTxF�
L3r��%T�;�i/��]rN&_�ǴP8[�hX�cn7�6������G��G�U�Zq���,�L��c-���Ǳ�u /���T�x��4����l�沈�}�N�=ж�N���(/�����{(0��:N���FWA�5t�D� ���£�Q��jS�����Ã,T� ��n�m[7
`{�rot�^jPԾT@"�2����8�DG���;? 컾�!��$�iԺ�Hq�6�m�ā��7-���w�3^<+�F�nG�S���'Z���u�L�w�����U3���>]��V1�u~	h"y��J
�b����꫻���_E�}پȞ��j���~��Ң�`Yy^w���-��.�g)-���A����>}�*�������W�I֘��191�;W�S����ɏ�2����u��b��N��p���h.��!O;i�ߞ�PW_��N0t��U?�%����&	h��6]<�)�#"w�'�Zha�&r�h`d*ue��L�m@�5`��no��z�ҁHޱ�����=왲Dȫ�)- �������c�l��s<����-�˛p�i� ����	��u\ިc@�(<��_;o8#	O�(\�5f\!D�G֭���*d��*��m�(���S���)���W�Γ�m��b�3k�(�S�eʠ�eo���-asPmF �&t*Gq�b@3���&����L���'��:
l0N��b�g<i&�k6{q�%��'��+*��0���*)�>9�`�>���s�}Ƽ|=LXzB�&vf(��7mG�5wȬ�x�6~q�7���w}��>@l��#{��$X�:eb�2ř-��T!g��n�FөA�=�έPyݺ����x�H�h�W	��ޒ�(��oC����8P2[a�޻k�%8�}���.���J����S<��(á  O�)�u s�̃CuG�U���fB.}>�: `��ţ�"p�^�ַ��.���Oɗ�g��t����ް�J8�(,�ފ5�lSӟ���<^�0���Bm�ST���#�v8��]~�^v�Ѯ�T��s'.����ˈ̵�i��N�'�.�	����yN�N���Ɓw3ꗺ�q�ǿ#�gܽ2McR����Sy���T�6ڭ�~#[鿸u?S�q�C�uB:�A���B�Ta�ՖA,��7l�5��![��}�KG\�앏�i���_6Y~E�a��{W#�Uϙ
H��ltȒ��1�R�t�����[����U��7Ӭ�T��/�Z�1
AX�T�u2�E9%�~ϛ�r����T.!oI�>��.��Z'B��0a��"�t��[��1�_'�MI�YO#qG��\�g)=�m=�r��K����bk�?,��N�]��ՋM7?���';5��v�'�(���_���Lr���,�V�ԽY�W�|\�G^�J�N���+V��
<�ĹON�&�,�gmg_A�=�#�n?���Jn|��M P�����z\�{<�>���I:�(Z���>�l�&<4�[u0+�1���&	��Ñ%�ȹ���aH��{����[��(����	��1�j��~�b�&
�=�����w�bq���~w[N���%_�C�j��MB�щ�?�T��^�M�\�$�����������I�w'�'P}!vZ|��V>H�1�4U4��V����Jp�u�nz���]���C�G��:����ʧ��+��]��z{	<>3����6�C�������;��{1����/ׅ�P�a�mi�e��ަ����M֔���{n��q�~Θ�m?"�A��s
���B5G��^�,�\?Ɔ�ۄ��n+F'�O��w��v{h8�7�t
T�Z��(��n#5�@l�5{#�����%a�cj����]·������H�+�߸�mo�xM7 �E���/�V7�V1�f:5=�
J�	�ܯ)�T��5��	D�Y�-�,P�e��T�P�
�z7e�טȤ9�6�]�j&zh�H��w�˂��DAҨ��ȑ(�hH@� ����p��%x���̺�wE�m�nL�%b  v?.b��͍X���t	'o��fju&-;>�J�,Q�ι�-��2����.q�$���Jj����gvΈ�O���	z��0��7w��|�pD��gT������.J1�F��% �
XU�@�A���ܘS���P�Lg�D���=H�J�K1a��˷�a�"v[o�/<�)~gQGT��cSWݩ[�<�c�
��t�i�-���-��b��Zo�t[m\`��������K��~r�L0.Jl�#w�bt@�`�	4âY[n ����|������qk�r��J1O��H<�ЊL��c��b��{2�v[�YEu��3���[����ܷ{u���ɩ1�Y]���\��y]Ų��nR!��M�Δ�h@�R��^.�\ZZ������#')԰<*���	�B*�hu��rV��#O
PQ��Xb�2�7��q�/#;�d`g'�8[l1D�(���Vt�'�P���{���p+��H���5�ϲ&�M�6��g�r3bb㿞Id�x��}�\�#sB�Fau�
�h#��Q��W��G�P�#C�Bx� p��i��}v�"�G�D㎚jdh��+GF���j�L2O3+��y̻�����
������� �=tw ��
H������)�!ݩ��%�!!�ݟ��{}g�l�k=+��dm�^�O�gZ�M�	ǷZ��E���4k��D�kb�4�y������Fo�	�x��Ji�}����d#*]�YRW�����Q�2+��.�5ۦ$�@GG�΋� ��6����w �s.d�����Q��|���
l��x�e�*J��1v<��"V�7����~9�ʒi�­���������O���x��C�s���;�x��:h�j��(��\)�?<���,��bٕ �%|��?�}��}v�jN�&E3ꜿ���%�L���~��K>��F�e
5�����;�#B6��U��b 7gq����R0YO��* o�r����t�#x�#��T��:l�4������G���6�3C��:V�?,��xVڈ�s��1�?���WΗ�TݬE�l��m�4V��~G_�z  �#�!,E�;������ �W���v+��3�_��#�P�r;��fŅ��l+ZȎ5�{�n{���e�s�̆�s�D�����Ҁ���]޽�����ϕ�;���"���MW;p8�RF�p`u�	�������.Q]�%��=�E'
��� M����w¯�qU�ɗ�����1
W%6eJ�w��˽�9�����x~k�K��k���]�n=|��/��T��'���43m�a��b[��R54m�_���w�gty���%Z�í)HS$�켈\���k�	)X�5���L����5�?���ש�'x�\���kpO����1�'Y��������*���=�-m�������(�\����?}H�~_�[sNC�و�����lbSr�Q��u�Z�G�=$/��~\}	���̜��+w]����ǔ�$�����L� 7iR[�m1��1i�Ձl��"�y ò�z���&;`٩��-�k7+_d�W�n-v�皤���P�ʑEi���T��OWc7Ʃ	�{<8�W<�C��,���@�-�����x�l����*���Jڇw[_ؿ�«�ʅ�'�<���;.<�X,�L{�5B�����E'�<����-�C� �L.MQ�Rzo�-�%�����P7:;(���ݝR �g�K00�,�L�, �����&U�|*-h�*�wv�!����R�>i�-d3甞�6���c���s1X�ߜ���Q@�T�W�iw�9*y/w���5�
ɭ�$�����}�u�l�4�k����uV^��! �\ ����BvS��*�ݧ��Y�4��R��U�w�5��l�����?�}$�~�+!T���ɳ�d%&\����N��1v#"� �m;=�.���A���d��oG��^�BZp?w�U���p{��?��#Rs��EuّGk�w��K{��g�za�B������{!ėﳫݚ��Lj~lr�룃����e���9"�V���=��t�{;�ˀ%�}���q̧�X�p���(���öp�O�֨���a\wTP�teVx��G�p�I~'v㽓W�'%Gt�VZe�۱ ;�Ƞ����(�MM�R2��W� ��x)_�%�~�����p�[�������ǧ�o�*K�O�B�ҼT�+hK�*}�v����l5��n��ے�0^�l��haZ3��D����X�먐Qz��|��;=�ϹkQ�,m��h`���\����S�opg������NH�uXp0F��p�T	v��eJ����8�]�Ӧ���X�po�@zx��{�|ىG��p*T-�h߽�wx0�1��ZZ�9�=ta����3W*��2����̯�)������;�>/��x�[���,��Rx|��3X��g*�k��'嬄��N�K��� {���}�s�ʱq�� ��":LSx#��f��yђc����[=�څ����g�r�ƞ�_���D4�feƚ���s����-τ�l��S�l�`~��
��Z���HR�ov������Ë�_���n�!IY���mz��Ô�7�dWޟ��)n��t��0����G,	c�uR&'��:��?wӼ��y����j�o�L��c.B�h��-ݮ�kz��V|*��,�r�=�D����2�;s<+�-lm��E�'�V5JIK���^�u������}�7`��p��bh���?�^�_dl����\�&���r(�ś�>�%0.劺Hq̞Ƭ�ro�$�ڿ�hml��L1�kXa���9<���I�2oxިo9��5v�����99��Lz��_ĕ��ޝ�Ԑ� MU�߾�O:$�Q�L�1W�V���ܸ��I�4%YO�*�៤�h&'��./�%�;��O�8�3,��/����sԼ�A��=��X�u��=	 BB����9?�+���4/I��'�=��ML�Ђ.N��|���Ҋūc�ɾ��|˰j�a=3veE� >�X�%	����L���]�,�l�rv���N|EZ��F��x���
-���,.S:.���&'峣��5���K���X-,V8���|҄BM���D|�ڌ�HR���Z���͔���"v���������kS-�l�LK��B���&�Z�����w�&����[D�k?�2o�v駈�A�х�}"�mR�$��)�\��ק��F"�n����)�)"6�$g݊�Js���P9�J�0�+�M����^���ev_I� ��[��c
jeLJ��+V��k�]"�PM�����dǂ�e�PA�%7b���-�e��Q���+����j����r܁�d�_�V��r������I�u�*��X'VȊ?�D9�W/^�u�w=�o�i/S��uF����l_�m}}Etui��++�55�q�V��y�7���/ݏ�,�b����rx�dc>�����U�n�VNե�x��
�����"�@8���y���v���+��%�ްa�.��n����ۓ�����ܿ�%�#���t�����O\<F�KJ5�F��~�N�&��_^��VL�/�\Ϝp�h��'�ڪxqK9��@��&�ڛ̂�f��c����X�B~. M��3��~��\�b�Fe��C�ָ�V +�V|\A^}�\n8'�Mx<���qZb�w�'2	`�=���Zh()1C���^����+�9��Y���4��J���{?�4+q�y�^r�Y0�a��sh�,6׆'�!�e5�CL�������*���!>s���ݻ�y�Q�XV�%,2i�i�"�y{�{[�6T�O�z2'\����J|X� 2۔dÕ@ 5���m+У���*g��킅�ϑ���kI�`a�
 m'Ts  �+E�/S�����"0Ɲ�r�������ą�Տ��Q�H����z�- �R��N����-펥������$�^�ޘ����Y�Y��e����g��E%>�a&1�ϵ]��y�ZI<KB��娞g�Xe�l�![Ā��rə�NG��_X0�( eeg��~������������uv�aoHe	h�^(���EtL��J��j���O���MXu����=�%��=�Gf�Q�~n��WH,V8�\�E�<.汕)��SG��$����9��:Ob�_��.����'��V��Q�����DB��`VUMM� b�qL��S=�pۿ�6���*�?9��\K�l��q�-^��2:0��RRx�R�}�\8�!�Py���i���S@��K�UE$�B�ٚ�/8*Zh?��#|�D�V�\�����ǆl�PJ!_/~��.�&��A�d�lQ���K��o��1�N�"ō0�R�H�K~?c�ʆ\����i5�C�0~F�eLT�1.�S���] ;`��R;q�`�A����Q�Ȥ�x��2�X�A��W����筭����o��e�]�CZ�	U�2cV���k��lt�^�m�]�jH?|�峊� ,�n^�T�Ϸ���_;�d+"7��<�������ِmYӯQ��q�@!��JS<)�H�2������g$pTA�;UQI�1,��x�l���"���/�-y���H�}v}4��`�����_�D�Z�ާ�d�U�+M��;d F���𛯘�J��IMƝ���W��!R��Nh!��0��ҵ�斋����qoh�����ٟ燫e���@�������T;����s���B��
�f��D�ρ���쫂�_q�?����"��e�C�	����?qp��z�O>�q�|�S�V��t��(���THad0�M#�v6ba�~���HKd�3�m~yvJ�;��H�V$H�yP3��g�1��+:��N[�������>�s�3��80[q���Y}�9s����{�ڤ��e�&�^6���Cq�1��E����hE����ߚm��e��<���q[d���&3�Z�8�i�C�P�����ɗ��J�?�6)6щ{��C����# v�W9m���J���}v'��!D���Ԏ��<��^w1�K)�AL?p��\�[\|U£����8YmaVU�Ta:�9���Q�L9�L���Ƌ���d>RLT�!�	�udc��]�L<�~oR�X��������J���F�nW��81�
F�����&="�����d��eG�;:�Д����
�ۡ��MZu��D�� z���C��.Fe}����0���˕�},��3ְ�M����ƛ�ì���ǵ<��%^�c�5P�����D��)��WHrp����o���ed���0Ƽr�Z5�נ�.�\N�Ф�.��^&���k�^�k\v��	ϣ'����t#��3._����9pD��`-��EGх��8��zK�5	��; "4H��[ы�u�,b�mnY�['�z;t�Ƣ�� ,��鈱P(��8���ky^�i��'��M>�dc�Ea��=��q_v�XVNIlQX4�y8{�8�Bc!l���r\9Z�mt?{Ν�$y������Q�/���ϼb�,y��n.��H����cIL���ܭ��ڏ�����HF��2%�S�q�����Uv�$>ؑ����gS��e��ļ<#��D,Lv�Ub
����_�fYZrohw?3�C�f�,O��=i��|�e������-Wi�.? ��A�X2�˙�����|�i���	�ScHV��a!{\1/D�r��R}`��3 eQ4m�HA3ߚ����z��/q�g��;�mH��c�`�9I�n���N���ʕq�9�?z\|p�ؒNx�F��!��Q�RNv+�x#3}��p���jeWÆsF��7R:-6�ص��p�2C��ٳ��X�펷�@�  ȃr��"����w�m� |$��3�ֆ��+�Pť�'������a=�.��
���E�1&��?��&,RU`56����RΐD�\�:�LM��}Q>\�.�"݈�
��DWj������&��7v&������b܉=*�@��
>���!�m���ې��K�s���ʪ�F��ǒ2��T��T|�8����P0m�% ɚu^)�c���L����
�I��Ju���SТ D^�b��\mj�ø,�s�n�>�xP���Ó�D��(N�w�Aw�3bX�D�`�����/�b���^N����� �u׬#�)�ȭH��r��LCF�2�]5]�w�|�eFD�d��zɋ���j��[\�����eeJ�+��q�5�h՚r迷��=����XK4a��^*���������ϯ�q�6�e������tmt:�ES����SƏ����E��qݛP�į������`�����h����8��Z+�/�Ǒ�c�G̼�u`�#���r7W�ט:(���w�&C�P䊎�Lr����|S��"��kg��}�`���T�S��FN�|�f�&�t��)��b/o)��,�k�����U�<��}&�4r~��� �v�t�E+Hs��"���sO��0�����LZ��2�K��^-��@��?&'H�pb&L�3�</a8i{r?�=��#?>D�HQ�^��Ķ������]D�.B��_^6xL�,B�K��6�&�X�Nj���MFĖ��d�Ph���-����E�#X�%�������mQOeGƽ�"nS�a�`�c��ZJ�������ָj� a)���!�lg���K�b����a��G�^.e�J��er�sa$�3�����h�����,�Ŋ�$�"��U��m��V5�J�a�ڎ@�	�j8%�*A�y|4�l����v���N��
a�j�Z�裷�/�եSBu&�䑑�Cג�׳ֻ�N��F���<6�ҽX�d�O����_-n���2�X�aکp�褣MP�h�\�ŭ�
�3`;8���)QkKF��aAҵ#?���Cp��n�>Q��#i�/���-��&�w��Z�źɹI6ԕ�p��������["�c���Ś����ee��ePQ6}����g�%9&� �d&ƣ�f���_N!K�u�����_;�A�M�}�!���a�p ������_i}�F�eUP�͕,�`��ז��+�7��HS����Y]�^w�c³r�Md��|��p��k��ts�O����_q��:{���j��p���5��>$ۏ�#�1A���b����@�1��眲0��-X�C��n�e�˕E���>�(�R��`�Î�����$��v� �����;Mr��r�~`9����66\��>Z�j�"�xTShf��Ը ɇ��T��P�Zb�aUp��Ft�S��`+�5���K T�ͥ�%I9���X~)\�_T�]?�4�<h9n�s�ʠ7]��~vJ<��n��l���������`ظ�zS{�(5su��L�_�s��
�o�l��<��q+p�f:���������߲Ov��\J}����O[J��O�����_�/�ּ�(���C�Şd<�a�!���%�W�* �K���]!&U�t����m��lo���+m����]�f���?Ľ.��6|^��U�����I�����Tc�TO��F�8�*�x����W}�P�U�'��}]SR.e�S��Kk&�+�e%��Tk��dk�)*�T�348tw���GB���5}��+�FFF|�v��ӵ��E�~�H�E���d�pٗ�9+���ŅI�E� ��B��~��s�����Ibw�&��r���u��F�!>���gU���\���=y�	p�k]/�i}οJ?>��� �0��뚐�p�z�M:��)�6:}�t�In�ߘ�{y9SM���Q���._m�K�dP%�M^���$�-q�Ǌ���ɡkR���G�$k#�8�>#�Dђ�D�H}u�D���̟�b����]Ǒ�5�d�Ub]�13"8���?��K^*�=�4&&�Ya����j��O\�ɡ=�6>	�=M� ⏸�������������ou��Sn'�.�}�Xa`2���%��7�#G�hձ���5�lB�&v��ؕ�d]>/�KH@�a�ݧ1�.�ٗ/��+K�$|�?�%^C���Aae��h�)�����F{�ʒ�����ż-������������=xE9�M�( ��bo�@�,<��(PM̥�������fǯ[��_A�|�3����6�t}�?����"DgE|�_���á煇F��
�N��'JG�����W��������"�\�`�k�l��q��Ф�D�E��p��Y�m��6C��Ќ2`���c�~�UY(^%���nv`����y0���Ǉ ~{=+O�s��j�Md ���H{�HǷ-Xi��@���9���"|5b�+07���UxD���:�wW,(��GX2*�?~<$Tt��b�ߚV��N�V%��{܊����4�=#1�Be������F`��-O7�˫<�yϐ��s�
 L�D�z��N�\�63H!���+��A�ʕ��4�M��3|����WW�bC�1���!y X̂IO6��%DW�cHK�8R�x�����P"u(0�������?����̰�bJ���(���CX�������Q��|t�$�-�n�W�Ӥ9��,���i���Sb׉1�&��'�"+� h��{3��x��s	am�O�̓ZEp'+p��� GD�?��@{[�A�@�=%�G��oM��/	����j.8S���G�)���/3��`���,n�q�x����h"k���x���/(1�K[�ٚ���rf��X��*��`���@<�j#�_w
I� k��00��T�=�$Vf�h>76z�H��%3���/�>WW �{�"��7k�
�Ys�� �ޅ�� L)%�8�� �CU�J�CJ�<k>/,�D���M���XQ��"��G�󞁐j �Zr}�\{$�L�Q0ܰxP 6�Z�l1��|��`^�H��E��HYZ.�'���濴����gk��n�h���`Ï��ߊ��r��G�m�}z�+���<c��a�||�dDt�LTU48;·��@���)e�7fw�}��p�G&�k�g� ������G�ݣ]e�i?C�C2��G�����=�^�t1�
����݌���4�w��Lnx��1%J�v��R��i[��q'���T]������P!'�_[Q��=?�ⰇO`�%�	!l���Y<sRۄ�<�5��y��o�:P;_p�T���-t�ηķ�}��,�S��6����0ڗ2��>�]8�뗡���L�`��xN*�i��nB���0��Үca�G�-:\�[�{.��b�M��f���h�@;�}���$���*���SK���z��ڰd���`�	9[A��hf� S���Ǚt�C^*���Nq� �b� �9񪨞�����w����$�ix؟-��:�j&�tQ�ǉ��[�5O�^����Q蹽}pOE4Ձl��1ǔ���@���p�q�*ئZ����.Ş����*�šA�=6 �J3�s��Hv�����5?&_�]��@��{�r2��M����4�9����G�$٣Ccv��1���(,�'� {����!-OQ1��c, �Q��[�3����_Ž[��-:�!.�6�/3'�H�[�=<�uU�(��^ꈧ�Kk�>vǿ�������H۪��ɔ�!T���w���f�)�,�孙����'\H�����E�m�>�H�rO<(�� �E�g&e��9�h����N��q�μ�-cL��֯��t>4��ik7��'yH��ik��]I�\S˻��_V�&X�$b%Hɣ}�DGDP���y|�&���G���B��u�q\���+�Q	�7/'�I��b�]+;Q#�$Od�,�
U����w�P���$i�3������Tp�P�?�
:���s<ï���95�b���4�]�@�����=��E'�9NL�:��~�@�L�+�`o<���2-�4�w�M{ׄv�#�v�AK�3����w��Y�B�L}^n2�Ɔ�̤D�� ;r
ۀ��������h��E#H��3��S�;����C���9Z���ĵ._!� ��::��i� L�mc�d5H���;8�g��vĠp?�6y�\�<r4�jP�������#��<蜩�'z��9L�<9�:�fB�����?y�lF)��������8}ZHx�/��O}O���``3�u���mm7��V)��Fp�����xs�C�+l� K��l� �D|'�� �gf����""#����̇��Tb��#�ʖ^a0���Ш�t�Xz'>f}�5�TQ�;dA��+�������m��va�V�é������ػ��QtӮh}���, �+*���3����FC80&��oй�e�ڟva9YQs�a ���۬T���(�{�u�=�H?:�9�z�d�,�ro�v&����������:Wލn�Ϸ�z�� ��,&��������@�(j�6Qx�Vy*1"x.ˌ���i}4C(`#e��u��1�&���˓���y�s��8��\3�~~��<��j�7;���d\/������MΥ��Z��8!�����:ѱ@
����H��9��X�沽𦑵���,7����(
��Ӿ=�l]�/��av��T�H�J�y[�T�&�?��A�3[�:��JA/w��P�a�)a�¸�B�TOQQQ%y⽅)vVV�;�`,�8N��*��?hH��)�ƌ��q߁&W=(ߍo� pH�T��=���G�uN�J`̃gd����wQ��L�S[�-[z{b��?�B��`m�$��K�X ����c�#&G�e��t��}d 4��&t����#PQ�����P�Cz3�;{D�e0�<r%�Ԋ�]EҊ�(5pء9��;5cڬ~���J��xh�V��i�3��j��j�$��<�� 3��_�}8�6�7��A�D�x���^v���a�V"d[�P���n�5�UY�U�S	��}G���+�'H��i������f&6Kt�ܸ��w7�^�)�W��d�y����v`lJ�H+�����M%����c쁘,?��^X��B�@�휭@�Q���|���{oX�9�Tޛ#�K������<��J�����)�
�=m�N(*iD �I�z�/f�	t������k��}7�Ca��b���(�_H.���	�����܈� ��F�gS�����%�����0S�Y�M<-a	Z�p �C��ȤD��5�v�w�B�Z4��X�a�Ą�%��
���H�K��5 8ʂ�љs�0�2B��߹&ku�$�V��,娋Q�� ��y�e���

��!���x�]�HN��ǹ2b��ص�VNQ;8�'�R<�7��:�6p�����qe£� �Ԩ<me|�W�0��|8�v[L���"�?)�r:�y���<qc����$�e���]��Q_.��
L\'�"�)!B7�߫���k�V�Vt�O"���q�:�ܞ��R���� �'���z0(�֎�v�C����x��#�>s�$�G��a�Fz�)�N���&*���w�_��`�/|C�qw�w���Wg�2��Y. mTm��h��ʹ�`w�O���"P?�X4h{A��v*�0�R���s����v����%�o���lI<�H_(R���[��዇�$�G��c��y<�@��#��v�%�6	�}�<ϊ������
�zƥ��x/�Q��|�8��w�E�cY9
*45by�"O��c��wU��fr�i�<3�rZk�98�1uD.ҾHP3���*�5��0��B�սaƹ�ri!���٫u������P�1�ա���"��D�v���z͉���jm����I�ǕH��E�r�F8�����.��Vw�8�7�>S��_(�R���J�������E7�<l��	��F2G6xR�-�<�`��`̡� �	f|Ͳ6�I�r^��'!N�z<x���<U�\���đ�^
d�(用�:��%�*�f58�}���L��OϚ�BR���p^R�U"^&O�����V�OO�c���!}�G����0v8<�"�M��DU���PH���M�9��]����rN�Zd�4#FB���,�~ʢ)�����6x1�y*kJs�.����ԇ�Q"P��<�壅�c�9�9T�����A:fm��l$���C�&2��8����՝��P�"�f0/�NF�����.���K @�g4�D����+�%�p���V�ٻ
�Ә�v~n��͈6H+tg�ȉ��=����D*T��ޑߞ��^�,YM��L��mVQE�D ]$�K}��ݪ���B��s���}u�#$�����7kH'y\��v����}@����;�r��K��	��J���f��ƦP�.7e��#� 3�R�b��Wfj��=�L)����Tڷ�A"����'�r��0"��Tc�Ļ T�%�(�w
�Q�4��GI�藢��L�m �D���O�p`�@�	��t�,�ǚ�y���e�A�#9��唉��v���)���r��"���ݭ��O�<�S2#ET�[�H��4#��٩*����0�y��Ep,��G�i���K���y��(��X�^�D1�s�0/�+��r�1�TgcI�#Lr5w;�+�v8}c-)}c��;�"h j��DF�0����3g�7w�7�lnQ*QH��V�s}qm�w��>sc��4�Z�[���w���W)�@���5�
7�~��bX�Tg�E+��e��[�^�	�=�jjl���L�KƧh �o��+FY^���lQ��'�>M���c�(ZG���Y|��SD����m��C�rId3��ד%bj�����񷽟�29�
�O��0��\���(��}�H�I��$e[���hne2��@p��n5�1�+H/?��� �sS���M�y40�iA����c��j��� 74��#*��,(J���ᶐ�u�������CulVl�%�P wYb�����uZ��ṭxo'�ި����Ó�1��۹!���%��B|+�;J˜��8z�7X
��t��Gx�e�M-yx��|� �l� +�v1��|'������W)j+`�h����fG}�v$�L�)i�@k��e}N�m�:5���~��y��h'�!3Y]�D��/]Ry1��]�&���ˏ�Vk��]S�K��˝Ȟ�c�_ IJ`�3 ��9���KU-��_��Y��=IetG5���@\Q$p+�l��:ɷYR�5¢��	O`��1M�W��ID�m���se�B��Ud� �B۸�ʌo��N%����$�`���o3 z�G,zZ��?�����t�/U����o�EF�������6��#�	R��[vf�oAwn���Z��M�c��4��q`�сc19Ka]��-M�<�$����:|.�RU�"���� �QH3���+�#On�I-�;�N���ɬ��;��K��B:�K1�&6���`�'������Yu�b��P�.�@��@�$����A���q��<	���M�у�E�ܟǪ�I�nG��ܧ�M�*8U�#��Jn8��P]�a>Wg������m�����������}�T�<�!E1�9�,�����m0󿞵V���7�h���*P}+7D�Xy��fȩ~#���g]q��\��$4��� �j�0}�ڗ~�(�ޭd�h���`�Jlu\�w���4+�_@�<�.|-7�'�*�y0CG�b؀"�I�D���p(�E1��	�X�����IU����H�z�z����*?@a �S�5
�3A'A��-���k�w ������)���«�)����D��2L�H�FWl	�& ��͒nR�LEjQ���4��M!4�6
�XWg_����U*�6@��׵�;^t�=7�g��[}>��5�<� 3Ά����U��[������^�������Wf`*��W5�2G�A�^HO{�.�B���YIL�ӹ0@��:���ׄ��թ~��z5eFz:M�=�7�.,F�L^1!�f��).s]�-懫 �~��줊���w���-ަ݁�g�����G�F��>;��).߿1K��<���@0L�;��� ��<(\3
m�׉�	�[�hXx�S�v�E!9/oŒl�-+�a���ʕ�,z�bOIh�<�aȁM8NXj�Yr���@��7�$n����i�[��4�?�8qM_{�<rI���o��mP�ؗ�q �R�0؟���cZ$0 �u6A����!�*\lL�\P��re�p% �Ɖ��T y�l��D��t���Th�KC���z4'nu0G�:�o�����Wl�-kό*��]�G��>d.՛"����&���ǵ,�o�o�����Fz��m�Rg��vF�XWʩ�rk�c:E"Х(���I�DfԷ�3��tS�{��} ���1;�bDK\ep��^osz7P�!n�;:�J(�f'B�� �Q�.����_�tI���pחM��=�M�Ų�"ޝR���tI�g���;�8����N+pp����*��R�.����Q��l�v�Gڑo�zK�W��Oĭ�}���0.>{Xn1
�,����2H�=0�����q�E�:���� �����r���=��QK>��ڱ0�Y��u��o��������	r����ui ��_�B�L�,Yb�BC8�vh8��=0T�ɨ��]3z�sq����r|_=�6ᇾ�q�V���'��[�:���A�ޜ%�� "{"�h8��G�A�2\��[�|xA�v�M}�l���.�r97�m��X-�{,���s�t�ԣ:/[%�wg���n�۵�0�4��v	�M�j_��a�1������i��΋l�jc��!�T��(��I&Q檼�?��-Um����@k�"/�ئ�+�ˣv�1����3GBi's���N���Ud�]8F-__#jܽ��������]Ty?����g;cp_����"�wBώ��_�҈]vX�Z��{��)kF}ȍ?"}����U���Պֱ�Wi��W��|�ܜu��;F���f�btw���f ������a�	�"��yF´��z݉(���}p��O!���j٬���2�`A�A�nB�*��}���C�C�Z<(p�TŦ��l�88|UΩ��ƙ .����CM��#��3��f2�&�t�<D[ �@[��.Z<�/��|wҵ]8mS��r�2E3���,��,���΁ظ��g"�VAj�cKM��_tF�T>!��>�N�>58��)�ͽ��ldp��XŢ�HC<K�S��=��j���[�,�A˲S<��Sz�=Q���� ���(�J �$�����?��w�*�(�0s �a]����"�r��I�g��Z˅V�ť{���Mq�/�r��)M7����>�95U�P�����4��ã�^�w�Y��nx3Jщc�������N�ĳ^v�b��1�mc�Avv.���D�1�z�on��D��+�6�/�)y9�T�n�3�Z1G����L�`%�h�J�m({ҫ��ĕ�>)�&�(r��	�󑀰�ZqV��|�%ٺ�� ة�!(]�m���|����b�\D}�1	:�p���\��vل˥ӇIJxF�4�C��΋5�z��ݐ����a�n#R�A�e�9	^�Y���r�I�N�����'��g�(�j��pY]x0��YpU�'/���L�Oȥl��Q?�nsF�$I�
/2�9|�d)�Rl�2����q�a�����t��Iz���dG�\o�e�$���s�4�G�1��T��*�q��$�����	������i��A��L�����%h?׼���l1�1|q(X�^��d�DA�=�%��JS���U\���*= $����S<��6']fkj�J�
!�3 `n�y��l�Q=�}�'ׯ��Xͳ�p�n,�aX��#D��p!=�a��M�r���RϰF�|x�랱��ԭq 2i	�p�f��@�|���t>h�j�'.�$�4(w h�n8Sl����4h���j�rf��� �%%'e�ڃ�'#PLp�z�����nub����s��RY��$�K@�]ބ�V��̸�*L���uu��38��Y��|ZV읥�B%-��� B�/Bi�`�����?w�Hx�h�{�@ԬD������`w�P�Z���m)j�%������ḟu�q����4Ӏn���&Q��l�F��x����ݗR��������#s�б��~+�; F���k�woԟ�/��аPD(՛�~��`kl���TH+�ʝ���G��U]3�9��c����åtH5�ZW
Er�k.&j����
C  r��U�3�����2�%J��2��?y�zE��_-]Y���β�nm�d #]�Zr@���H������(u���z�>uWd4���+�q5�4U�_X{��Z��C!����;? �7�A��%�j����G�Tf��� Z	�s2�񖸩�vQ%N�Ԁop�����Z7c
zDR���WY�\x�6�������9���4�r%K,��B%!ސ��xA���@z�Gu`�����Xݖ%ĭC�}N�^�߱*g������Y�転�p��n�'K�m�]�� 5k�f@}�P����"�ܗ2�3����V������
�u�j�,��yv�M\-a=G��*���5G2�HZ)�N���2҃"�y�*��� p�ɲ��r�2��m�pȦ�B~�L�Pr҂L�w�i�\՜kf?��Ns�-��o �q���b��+��`�踔��N�yq,'���!�w�=r��׬����A��2�� HK�F!��_�ysV��#.5	��Ӽ�,7{]��V��
:�c!��t�.e̎����/!e`�Wl �n��t�5>^�'&3��Q�G���U�����,����h� ��	�P(\�K
ŝ-��8�	n�)�š�k��C����;����ޛ?`f�{����gf�A�~�E�ɪV0�#�LD�Zp(�x)�G���D����/+9K�O}CJ��B�Q׺Z���,�D��5���G��{`|-&,|Q�)P�?�}s#��8��X֛��0扨�nHS/S�V,~���]�ć�xj3��^�M뽼�Ռ�Z�����g�+����c a�@��D��l�RS�k�\���� C�5)~�z���~�$��	n<Gl-J�}"cUB��"Nb��hc���m4�� �ߤ��!s���g�*�N³�S���^��B���U��
�݃�a���?u(A��6�3�=z�M�&� 2?����L�F,F1��@	W�_}l��B %Z���q�x���:;i��ڲj%��Y��EIW�h���q�Ed=O�����,���z�(�,�p�L%��g�ڸp;.M�&��v�4�QPfN��}���tf��*�����$�7uթ ��6�p�c�a�`�M����~m�oN��r�ZRг�ii��oӁw����7a	�6�	DC�|Z�ݛ�Un���x��3��[�>��u�N1kJ�ht^�D�pK��C"����,�|ay��. �q�r��A�V:�i�g���:`(�X���M~�sр��Sʔ�Z���Sg�B掍@_�6DZ�)����_�G>�0��+v]�(�n�=�6��`O<f�'�,�ℜɤ�( X�@��9
������}Ъ��L���DF��8'16N���C3,���UXf<��,�2g<���p�_���F�u�w,��x�7�r�cB-'�QQ���ӗh���/D鮗�g9�����þ�I��K� D��͙�	w%�]$�o��k��-|G�3'�㢵��_�3�\yE�zʳF�pp���������z�±r�UeK7ÏqZ��OV8���ڃ@���0<aխ�O^=���Om�dlsJ�C#�."ͼ9�_���E< r��u�D���+�A�'uU �Aѥj7�=J��nb��Y��u��|�����O�+K�Qi���؁��z,��~_���3I_��GV���[B�?T��ҍ�x鞲�ͯ��D����<��3K�l6nJ�m.��Ŏ��mw� П��7}]'*#�/P��})�-�?�0�]��{��	AO$.�2�w�$�x'�+<��y�:��C�O/Cv�n�n�.�5����!*�*�7F�4�2#(�/1+�6�Ц�	�t�>Uff����؋#:q#�N|��̀�A��F�ɏ0�����I���{q�����r���=/��n����9�X��/����]낸�����s͈�t#��o�
Ք(J��,^d��Y���k�1?'�Pv�z�m,���'��Q�z�v�j	��{\a��,f'��䤉9v�9�i&!���Q2��Y�G.���׽�P�݈��ʺ����6�9���������i���-`�Õ@�gv�V��8	�`7��)����g�!�.������,�]G<�l�W�A�C����#�\�g ����؝pq@��3��6����˹��n�7aFF���L����[�%e8�g@00l��l7�b H��bh҃���Cf��9�����&QU�p��n���|ؕ_T)c�R#��j�a���_1atOl�`��u�N/�	����4�>�yi5f�d�����~�'�(U��\ z/k�.�wAN�U��Qe���*��ZI�ڄG�z�&����Z��Vo�;��tП���1Яv��f���T�B3����W;s[��cʔ8�99ӵ�vCeV�B��3���G>L�Z�W�A��Y1v66��%~�cU 25%�����8;�;���;��-�k/ɢ���t��.@���Ϙ1��&F��K���q}��]4�o��HO� u���݋8w��.a��$�w�Ȅ�6�7�Qϯ�	��͐�|<4	~a�~		��~�gc��4Nu������v�:3O�#m��ezF`��?S��G��kH;5\5|9g:ߋ�s��P�K�gQ���q@�+4JY�X��@�5n��q�����I��r���㋰��|�8��L�N[�������¦�OH�
Gv�-'X0p�G�Ԯ��|��`l�K�y	����$uu+D���~�h�ڬ���ξ�b]����\8��`��,s�])5�E�q;Mlr��i����H#�F����FoIL,�]�K��`�+��ߣ��#�.��³~��)��V�T�)�����7TVMnڼ�φ�L�� �y" ����7��VǑUn8`7y�WO�Sl�re"\<S�\�P��*�aB�=�w��l 8�e �O>�1������{&uE�~]��U5=�IjX�W�/ΐ ڐ �	�|����F��=���]��$��`0Dp��Q�:�����Y����#�n��Kwi��e����6B���ɣ)H�@����.|��+*�,숑�Gl���h����9=j0C£^����U����z�i��P���6 �ɚǷ4�Xju�Y9�E�r�U(�8ȃ;�ii�i�Ĺ?z�o!Z���t�_�
?�ː]�I�E�o�2O�qW�����Dh�	?=/}GJ�ڥ���FR\+˵'G�ix�M?T����f+�B]J�R�*A7p�]���c���Q��=;J@� 3 $����On:���KBJ���$q)g!��D�|�#��v&���9f��}�+���{�rM�/^1�\8��f�_W�� �W(�̧���bY	*W�����&���>+���}CQ�ï�1�Z�J�����	��w2�:� p[��?h�TOy�+��y�Tm2�j��ch/s�� �䇟��Vc8��*̷�٧�(^W	��B��&�U��tUUJ�pl��<�.*��F���0M�Ȱ�J߻�~�5N��v��
�B#�Kba0@��9�=U��Y!���ُ��![ח4N�8J[�\�"��V�Rt��S�f��{���	S"�j�ʵ׶WO�@(.�אǺ H�
&�w��p�j{� �D�^H]L� �v�\I�Ѽ�&h�pݸ��e��z�����uD�ܯ�w�V�wQvN�� �< �H$g���V�W��Ɏ��8o�tq4_%��ߌÏ���a�-x��@L�U ��{��_/t���Ii偼���<���H���'=��X�K��=�bV�`~�ϧ�\��nu���Vqa�ᶕ��X�B�ؽ�+���J�67�y�X"�,%�K�c�c�;.m��$Q��o����H�&3�P#Cl�,V���T`�V����S�1�L���i�f"6A���0PLW
]��T�bH��^2�]	G�QRutqo	U/�B%i��A��TÔ2n���j!��th�ۛ_���h��11Ϙ�"�4��ޣ��̱tг�vd��)W���o�ŻV��k� �:EK�Cw�˽��IV�<�ԏٴZ�$v�k�cɆ�J�&2b�m>h�8���`1���t�'P$]N�E}%�W���d[�0�'!�Vb14ϟ|�>_�m�"�^-,;]/V��&(�%��A��X���
V�kI�����BK�W�2�gz�KH��n�!{M��
P�X|d�o]�
hS�x,�F�q��W�P��If�m�7Vo��o�j[K�=&
2�����[/���P4Î��|+�N��j�0C��*�2qe�?��W�v�;���vq8�'�����Bج�VU-$��ܼ�K��T��BAh�x��ZB� 4O����>���O8=R��4�~��(ZJ�H�`סݳ�ЅD��}q���{]�T�0��Y�&�j���lq����͢������-*]C�,�Bc����\r��,	N�C3r�	퉏z���Bz+Ƶ�LfDE$�X=�����7@Pa�_�d�3�M���1�'��s���n�	`���2/͟��d�GNNz���J{ҝ$�d�U�����g�HY�.  |L���-H@cJ<Ȏ���P0_/���v�0Az���㯀��_*�l�˖3�@J�6ɮ�G��^��N���ezI����TKnRً	QrW���������t�(���{�� �mha�)&������z^덵�Q26�:k��/�T�����^�bػ����c��߇������E�]������֙���nD��K�
>���)��3��v���9l����5���\��^��v��ѡ��]�Youb�� ��{8�\���T�dsv��'�i���C�\�X\L�9@ٱ����C9�9�� J)R��0T�;�40d`d���i��/<�W-5o4��5�R��٠:��m%�Ke��{��x��;	���t/��nW������1����A��2#�Cq'���qv�t|��S3�am���K�q��N~����pݛ�
O;����c�}������|�t�1��).~6���Y�i-�R���/:B;�E��->�Q#�A>l��D�6D9z�	��!p1�(��l?`r���S���������5K�m��GW��.�b �"?����j�t@P��ّ�+v+h$��MD�����j�$ ���Z���OVj�nº�t��s��&����v\<�sS�D�z���ǀ�m�e���w��}	[bN�1"t��,ɪ��v,���y�B�O�/e��r����0��~0�{{!��b{�������v����E?ϴ��>�A��_#;NV?77d\�Xw�6(�q~�A(���kw�`g�w͊����R�0"���|�ʁ�k
P�+`=w;���O�K�����'H[K�?�~�i�(4�������B��i��jP�g_�He�.s#t4����������,���y��8��G8c �R5�L�٭V�BH�"������#�%g7÷��H�i4m��f&�,+�b��΅ߢ-��d���]�
�m��Ʊ{����C��uX�*�{��Qf�'p�A���g4�N__J/�=���n
����J}�*�Aa/�h�\�L���Ó���a~���lވ�^_E��[,S0xͺ�-���%4��f��ᡢK'���{����ݩ���Ipp��_@r�خ|���a�/��ce��VoG���I�Ђ�{�L��SA�����3��x��TV�x��/~_c�>;�(^O��7  �0��GN~�T�ߘ�,�j�/�o����!����;���ux��*\(�'��� C����~��~�I'h]g[I�o��h��o"�����/i�԰�R�|����*G-�I�}m!S�i�yFP˗߫�˓ �;TCً��|�%���L�Ɇ���G|�m�wHN쵭���A�q�Q1"X���6-��\����"i�f{���!����p
��b�x�P����l�Mq��M��H��Ԙ1�h�-a�6Ry�[�tʫ,.��&�-^#΃�X�T�V˸�#���Q�U��'�����F�k�u:0O��e�z"�f{�b��7�F�����B��K/�0/m����jEOYE�W$��e\63CT '�����k�&�ͤmZ�䁼�L���k�?�1��������������2�T��������-�۱i��JI**��^��R8��2���=	�N7���x�G{��*{Ͽ񉍠/#�6��@����`�f�Ը��J�-�j��p$49����\��~B7��&��1�q�.�=�ɨ)����x�.d�%�0*����<�b��@�ev��ǍVaꝁ[��pΗ^p�Ο/D'؁����B� EzyJ<˃g- XU�:����U�Y�Ѣ0/b��g"���0��X	c� ix}8˙LW�$V����3Y^�`b�(ٟ�ܟ9-�e���V�t��� $�.-�E��O��˖��|���u"�H���B��M�Ж��_d;��**OD/�/OV��j�O�u��J�f6���D���[؛c:�5[�{��}��
��"rM�l����?iT�z�����[ߌ'_��Գ���p�싄4 !�B�MR����m�܊�R�?���N��H�i�,��,@��p*I��qYN"
l��f�)�(b�~ހ�#�Y��l�4��:ȆD�9��uqE�����?�$5ah�"�ն�#��вɠW@����L����Ԅ���]��F���৺�B�m\�"Ĭ�7��lX�ԋ�l�#�_����̂JsHp��Bi��	�zrY���,zu�\y��Yː��ww�@0S)�SJ��w3����E�~��d��ȣh6��m���b ��0�5m����\����%�銁��cѦޚt�y���U�u\��ma+�x�tw�U�$�;��"E�E�j�L�/P��G)��xL$O��!)k/D��P��O��H'I�����r;�J��)���>-d*����/-d'0��� �%5����j67���mjpG;��#9�xM�#�t��#�V���V@��9!
�����X�:���d��!�3�/�Y��v ��϶�8�π�z������� �KGl�F�2�h���5o#�I�TL�Q1i.tz�}Q�c2��/i�	j(u�h��z!�$�D��2�
 �i ���PVU�M#x��J��Pj�s&���GT ��*�q�Ю�b/��Nx����}Ьd(���Ę��f���Z���:Bϑ3O��VJ�:%�9�Yc��^��.��3��	�E峃x{�E>�pm�>H����̜�?R��X nM��J�^'jj��8Yi	�����8<����-O��BP#OK}1�����s���v�e?�1��oسwG���#����f�B�0�����>;�x�/�d�\a��8��k}�F(��:������ȷ�������N[ek�%<�ԕ�n�f��oD�՜M�v���f�9V铤q3M}Ψ��S�(EG(�DTx�3����sZ5�z���kcʏ錷[h�UG�����M�B��}�`O@ZE%��١����^R������dqwխ?��3w%j1�`�Rc���$��������!��Q`�%��b;*"O���
��@~.�Ŵ�sp���0Y��)|�$��� �4Z<Jd�8{�耋A�� ���-/E�L���<7�k��sZcV��21�o]ЩoAq��["�v�ٓ-%H���U~�xz;���!�"�67�oD�|s0su�R)C�W.}�����+)OmÓ�&�� ΁Ie2T�><S�)}ZJ�dC���P�Y��5���k*�J@uj�$}g4��KJ���A|���Kr�Ǭ�u[��DU�F��U|b��L�*�[�!%X�������})��qN�窒>�A�:��b�`j_��	��W[҈R1�'�dK�.�=B����9'ā��P�<5)5��g��?.3�!Z��j���z�J�5�:�ķ`}�����ʀ�V8�vyj����M�G{X(�[.��q�p�b��X��%ֱ0$&�ҝ��+��Տ�Y�kaF�8�tC�-I���3L����pZ���#Y�X�8�I�
�"z�x� Tm�6Ø�@.h�,C�'��B���鈼i[e
K����~�|��% �Q-3���&"|=�gYZf�݆%Wdza��( Q�
"iLdT�z�E�_�?�ٚr��ZJ�p���G���J*RX����xQ�LX/=��>8��~2��[ig%(t-7�Vڔ%��I�X>K��'����U�����ܹ!Ǖ��h�D	�]S6��EV��.�ܥ~�H	a�������V�Zn�z������כ5�q@�abD�>��:�j����E6W]��H44-utr��U���P�u`����]�t�](0�,᳡٦�=�.����	 ���MvD�lb�'�C/�ݛjjaU �!�`&�8/7,�eFE������o��p?f�����A����zE�m�p�˴���z8)=�;q���������EfO��f;]~��k;Nt�'g����Ӑ*�L߂�+IϺ���Ƭ�0~֤�D)�I�kML	h�@� �$��jt)]��Ŏ>�G=&�č¯�-�z�|+WYAY�:�WP�Ɇ\��#��k�;p�SWea�J�Ńa�]r�,D#CL��P/ޝ�L=���$���2{�L:�>|�A���5rhң��g�K�<E���s[ߘ;������Q�ý�����Cd;��c��r�(�4i�
9��%��U���Η��7�$O��9� ,��5\m`â
�Ő�	rk��������/��Sy\-����d��G_zP�t���w�g�o�X�x�1/����Y b���{8�/�.T�CWO�7T�%/��$J�-������&!���<�4�g�U��&�U� j=�#ή�=��8
��Q�� �~����ˤ X�[oF�"�|	Dh�^����~x�x@Cd��"�r�NK�����{:M-�X(/�H~�|���#,�N �="f[?{c�/�u�m<�Tʳ]���b��m9�c��H��6M�*o�O�*C��z�X&�D��(��r�2��V��̽�s�MNb����Nƹ��\M?��L�;Ia$�m%B�A`ǷC�ް����	�T1dS�����I{�]�"��-�գ<�y�)ț*2��fl���s�	��!�\��w��q.��0)7�w��e�Ko.�ʠ��E��J�J��!|x�MBu���p�h�����lw�0=�R���Ђ�L�w��h�[�����l���� ��F������K��z,ϟayޓ�%�dqf�f=]�l�z�S�&_6?ֈ+��9���Yΰ<= z}��'qx@3��r��-��l�br
���?m�r��C%�c�)�1f�I�?�Ǚ|k�q�.sT�$�>��+��{���h�Y�����Ӈ����9cd(T
{���(	o������N��bC�3�=rQ_��iHΝ�]�>�_�E��\iV�1KNl�&7�j��i�I6D2����g�O�ְ��}۫J�>���t� �c��n;�d�֏F��X^�Ř��m����ʜ���ZE.��k���M�:��ٔUy�_0]����_�IT$�h�~rΗj3�������W����*��#��d0���7��\R�Q����H0(�7�Ʌˉvv"���C�v��7�5�ԋNV�S�A��O��D��_m;��co�.-���wE�:k��m�!2��f�%/�[�4��jM����y���FAѬ���-�sR�WeR|E�G7����R_�pU1��@|62K2"W��Y��^
�Jq�>X������ݗՔ��[��n����R*"��V.��'�X��`�{��e+]����2H�XH����
���â�d��  �b�XP��	\�.���>7��,���Ռ��gǇN�{�"����T>S���d]�KR#�e���A�׻���c����<�׹'f�j	B�S��.gd�	�^H�^/e�Η[[���I�qZY$I��mR��#�kq�4�〾�l|Wt1אd�����ݭ�f����Ѷj�ｶ��Uk�?'x�c��a�c�EB��͊�2�ʊ�?�����h{3B1j��I���}f3Vm��C���ɦ8�-_��r{�R�i	8��Ͻ�R>�9а�j��;�"�ߺ3kxb�'y�ki�؊o��QC��.��DO$�[5�ySh����8

�����@M���-�u_����h�k^��7�k���Q�� 	C?����W����cɄRV!P
/ډb�*4'Nã�
�`a�ؔ�ct��S����O�Ej���\"z���H�R��>j1�v�`?��3ʚGǂ���Q4��xk�j��7�0]������#����
>f�\��B��
�:\�G:*��@~��D��㙑"�����X�厼�K��;o(+�-6,
�о��Ò�Uf��U=���~��F�#�q@'��H�/��T(����1��ˣRRsKJ��$zC��.�u�i�Ǩ�$�tk >6xh�i�E  �gEEV�%k��3�"� v	��|���祫)���m�L5�y����*�X���4N������;�@�'��kM0�����t��H�����;_p��ݗAt�r^1^n����qŲ�͑h1�O3C�w�Ub[��!�_�-N��ٱ>IJ[X�-h�s"��[�.�Fe��
��ku�c#R�g�p�N����3�_� S�d����q��5��]�i�$��GU�l�����D��'G��7*��Y�"*33��/�^�^�᥎�*V�S-N0sjT�}���XR�:����K��Ù���֣�[h����Lgߙ��79����r�P���Ԑ)� %�%��5�(�4��߽�E�)Q�%��N+��rI�dC�f�A�z�n��� �[�Љ�� ؀����ޱ�H�\�{~�6�!ߥ֦�����Q�Y�i�HC!��+�m��C�Ă��c �Ǥ����A��ߊY�kͯQ�4��T(�w�;�"��l?/����蕅�'�&�%-���*K�� �3XW'�o������g�����5)�g{�<y�pݵ��A�6'����O%.�aA���}a	������X�	��e����;�/�ԫ��K�f!^�ݶ�nt�kY?K/�:�d�����/S�t��c�
���]��!O�-�M�d�ݯ�MR�vLc��C������/BW��w=i���C�Ծhyr�+ �R.��:��t�N	��n�2�7D_&R� ���&&W%Ñ�	˶�
���z��0B�-����;:�fD���yz��Cgk�tP	�?_����	I�X��6���]j��1D��BEB1Fp\�r�o�o{�li�pw��� N ���+>Bm�:�;���Us�Rа�~�.)H�������~H
�>Z|�=J6�{{ g"[d�C>ZJ�V}��zL5^�Wq�}�����k8q'Ӫh����ޥ'OXߔ��}�[╶y�[�Ιׁ0��(��W�2^�qmcy%���ˊB�
�⩄I�O����Ub��Z�3�u����XcQ?�:�.E-~Gq$����$�>�l8�Ώ��!v������IMm��q �6���n�
�Q���t��ٟ�����r#��/������+�Q��҃�� �����-����t���_��/��;ש���ᅊ�M�ѧ�OX��E��&��D�<�o����N�3��֢kv��3R��&��W�N]!�1���`A-��E��r-3�����/�%P�����/ۑ�~C�>�b,�n\����1KG>,�,�ݒ�ES^�7���QQiHk}ս�W������@�U7�	�eX�>�j���bm �S��<�|���S�`�	<�%ě�)M��(}���xu$J����VO����ER)�����q+\q��@T���Ӫ�r�P7�����&uuN˅�7m�y�������U�Q���qB.����ܛ�o
meFΞ�������x��!u-�:j�1���H�Sٍ�A��5�(��/0���3imN�mB-�t�J�l}-���d��*G5]8
�\�_@�B3�h�tH~�A�R�jP�1h2����[� ��)��8%y�t�<)"床.L$�	�>���y9�>�#t�)D��v!.%� GX��Gn9�RZRn(*��V)����u^��<��T;�
����:��K5I���;���Y%�8d��Uˮ���Ex�	}��ː���Fyo�.���sǙ�����~eh-��b��B�4{yP}�wt^���o(��F�d'E��?�T~��-g�{v���\dE�u��r�Xc��J�&ټ�2�	D��X[���oQ�~M�lU{�q/՚:ԘvF|R�Wc�ԁA����q逕��q�A`�o�$כ�k�QȃFI�	�йGn�.·R�3�.S��I�F����Co[0���K��2���+*�>G���r�����I4=|�܌=E��?'a��_�K'zu��?D[�n��y��h�i��)��	m�L�º��2��p�%�Bze�;�8|���O�<	�G�e]H7-����N�I^��W�%�����;"�!�%��P͚�N��;�,*�(DJ̿�0�`0F��L���7%֕+ӧ+'8�?�A<�Da|p.����5"�9�{x&��S��=��J���hIJvL�'"��RZ�6
Ջ?mZ�0���r~ux�C�`�A��_��C��^��d'�F��m�4u�H�C'W"'�g<�_��l?Aܹ>��I���1��!��W��N����V��|��3�eF�'q=�q������(A��]^�IF���Pwaݼ�Y����z����B��!.)�u�=�9@����	)����ph3�찄5��?A��]Ӡ8�����	A�[?���3�%�����?��A�W���2�GZJ��]�,�Q|�;4{�bC�WG5�6䪶'i��+Z������S?��3�6dI���?o����^[7��O��B�j�M>)����b���<�m37P�0�{�5Tp��8 V�S�����e��¿�j�������<�h���p)n��3!�_����dK�1c�3�Ո�m)c7�Ǎ����e�\�\�0d�N޽�:�"��6pg��U�+��cm]j���46�Ϣ�/��꘏��Lߡ�.�s�U�E.U��򛽂}�8�3�j�!��Ld
.�Bx<Iɹ������CX)ƞN|��vhmU�^�k����F雇�ƾw:=[�0'��l�T�>�eBq��E	�zYl�����M*,ĝQ���_��HuЂG\�K���
MДkc�b�^�I�JSg`R�.Ӥ�F�R�M˲�Ì�����&ʣ������N������n��YXuO����3[z#^��s7ۥ
��#t���:��71婺�܍�X���dQ�W�ވ2����6?��+��uz����Xƿa���\ZO�~{8:uMS��������K}���G�M�;�a(.:���-3nWt��!���"�El�m|?�w�.R�:vRs�$�;-���yWI�!�"������z�w�ZI�N���"]Z$��p�N�pVd�`���F�G��ww�?�H�ڭ��#��TV���LY$��3�S�dsM�F�x�૰�a[ޏ���7�9"VT�U'��X��Jo�/����������p��������O�����/���y��=[[������7����d�9�s7� E~�?ܐ@[D���MrkP{��r�[���]v3Ja^�v���U\��'i�߫�|��/����[�c2E����3b�Tȁ�&߅����+��������;�xiK���ܟ�R���S��8I�n8,B���vŲ!).a+�xO'���̘��?]+�{�NGOR��Sl�`r#�����B�y�/z��J���,32��� ݭ(�Î?��k��dJ驇�]� �w�G�[�Ż�\���<���~���C�<�ԅ�rJup,z�0��,CY��{�Q�o��c��ihŋ�V_9�>�`K8�����L[�3�ΩP�Fn`��.{e��yN�d����J��!S!#H��6��y��oEq�q�*ܮ����Zŉ�ʗ�>�4Ŭ��,�7qlV̿}ݰ	q�v�g<�X~X�����}���ֽa��b[���:]z�!��w���b׶�|��5 �g:�E���Sw��@���ɪ�{k�V��V�����: ��*�o�K�Qk�6/w��m��V��`�4�,K�N�Dג	ϛ�=Jc"�)��M��"��w��戀����u��wթ�0����E�@ ӎ�D�Fv����Đ�R�E���ё���Ρ�&���1Z_���Ϳt����|T���b��?r6��M1]�|���M{�$8R��ˢ��ᜯa�%F;x{�{֗`Fk+7��Κv7|����W��^��6��|�ܦw�6�"�Vκ3��7�Ye�a�Xġ�6����"�C�W���tFe�~���9�"*ӽm9�b�(zҐ���9˃�7j�Oc:�֩*ej'��K@�MT��W�E�m�T�!͵f���L���k�����wV�wi$��Ds1��}q7��q*�%�Q�69.Zޭ?��90-�V�R�����J�ӜFA���J.d�G��QЗ�<=3�f�l٣9�(7.�Gn��a�2,��o�&$�ƪ6ǡ����ޤ|7�9���`Xx�W�L����c�~W^�fR�@|���u���b�Nx����K�b���X�co�=�����C]�<����W���ZQ�&n��q�:���	�%�~���$�Y5�ugD�+�����ț$�^T`� �K�r�����p���^�l��+��ݑ8�	����5,|B��Y��my�a°J�.���`��Gl!�����]��E��j�Ta��i\�����xH��n��xGg��OMWDhn:�ײgS��w���:W�ZMJ���b�����T&������5�M�éƮ�N�!�"�����P+�oa�R��%Bu��<{�ƅ��"�mX�T�&�*W:�TǱ��AH��FSL���p�}�>bk��AЌi��|��[?�o:�uGÏ�č5��R��6`��&D�ǩ��)�˲�-&9���u9i]��d��~6o.9�z�_��n������K��q�-�(ϭ��=�2��<��Q����K�
����-?�&<����B��1��u���6\��O�ʧ�1��:�de�f�A��q:~���o��9۰Ԧ��\��]5��,��f�oZ����5)Z~��a�iS����He\� ��o�آ��"iW��k}����}��Hb�%,�����OG�=�m�ʚ޽�,�Q*�:^K����s�ߖ����h�Fɠ��`�[�,��c�k���/\3�0�3�Ɠ�6��C<^#&Tf��ֻ\��Y�W�IvR�I� �����$��+K?���j��v,a�a�w�P��Y�~4�2@���ч�e���<Q����K?�$d��=J�f.��`�
ĥ矦��u��xڣc��7"Ce?��śm��'8�(��,g2�Si�(r12@}���P�q��1�n�A�$��M���͓�y�	��_'	L��Hq�<��?�Y�]k�͆�'��k�VW��	��+�f)�J��r�F��Xe&�k��q���z�޸��׺�`#���C�8���@K��.ov��O��?�	I���=�lh�L�MX5�\�l��&*�@M���I}�i^�"��j<��x��ξJ���"6bI�����k��_��D��2����T�:o��\��+.28(&��Q�� ��eN�wP�o?����j��W�30 �=v��R�J���)�)w4z�*To�w�O�i�-��Ep���[�B���v�^s.��
Vǿ���t���-��ߴ�&0��-wE2���N	s�2=K�
�/�ķ����\�Z=�+����ËO�Q���Aȁ��Z;�Wl�+������7F7�N��OMJo��~.���p��D|����j� ,ʼ�����z�%u��<�Z�˰��)�4����1��;rR�jgm�p������v�7�ܜh#��1Bu?�B�������DE�j�jZ-����C^��=TNeѪ�
:B3�Ajs@V�S2~�_:5u��B�¦�<f~��Wu������F}C2o��/ nx2�<�k��g���d�W�����[��y|[�}ʹ��"����at>
��Y���2%͢�����du�K.�Ű6Rd��q1���K����~�"����'?���W�.���C_�j<�I҂���(�9��Y�����ؑ��?:{W�5\���L��KE�n��c"пY,��6Y�]��u7ԭ9W2U"�u�\���Rf�}�Qm�d�$%��Q�RZQC�\RUO�wF��|C��5z;��m:��	��Y���/��d�Tq"q�Ǜ%�3,F-�U�T�2���+�f�y�^T�yip<mh���`���;m�r�0��~���٭�EY~���J15���-v)acS���K�7�j�'uxC�%8� ��ǈ���Frv�G���.4q�����vx��?�K�'=ٿ�u��SM��kNr��$�~��\�y�aU�m��STk!�<�/i/������]��PZ�DJ����ˋ��xyv��ͼa�'e�g��gm��m�	1�|{`�K	�ʔ[{�U��'��p�g���<�G�[?�ߚ���w�U��O^ ���>UE����ڙ��J�o,�.���_G�̪~&Eg�?,��mߵE2�z/f�W����e6d��x�y�~���P-�Wk�R�6� H��3_m;n�����?#R��j�,9 {:��hjh�m�����o�������"B�U������f�L�$y�28OөK��3Lf�'.�o�'����>���!��Y�L/���~�4w�R�u���o�ʄߓ�Χ��l"������[�|�4ɒ�@S#l
BFp�pH��.��S�U'�1�@h]�NUn����5��Nz/�n�C���/fu�c�cP���8���߰��r�V��R����@SM��x�%*�D �mv�m���h���c��ho�	�]�#\��Ff��15-�[��ghy�y�~���dI��]l�\��N�ѥ<���u����A�.��0]�eY�"J?%h�Q<����QH������{(~/��lI�֥ƥ�L���&�}�3 ��0�/�;'�u��lO㤶I�0N5�����_��"�%6����*�+/�j-C����Z�7[����'��[u���O�S�!#�����å/��}���0�JO�{�`���W�^�"%�? �V��Ry��-TҮ���U�����T|{c1��q@����]����.<�Y�P;�&
��ه�����?
}��2�:PUG�΢�O�q01p0X�G��k��>�ָ�Q�)�|��Ql�����	�ݫ'�b��Ҋ.��(E܄�"lY4��Y�ps���m�����	ho���[Uip]��'�m"d�C-m<^�I�c�`j��'�N]8��:�2���I��E���F�t~B��O���:z���+_�~�&����v甀��v�u�w����1�n���9��S�3s8m,�L\�©bŤ���ޫ��&dj��t!|���!ׯ[<�����[����$��L�b3�q�ZG��6��I=.�JLi�
Rp�4�v�	xP؟��^J�8�05� |�%�7�؞�����\p��FQ+��0��qv��y>`����!8+<��#�3��N͜�6���cG�.�F��8�I��Q��|��F#ۼY6��X�Q0��~m�.�ٜզ�4��wY�[�Ux�k<M\*8��9AM�c�ڹ�|kw�usվQی�y��lgM!���6�B�/���4�5�V�HǓ��"qhYٟ
�u�L���v�oy��w�gǵeUnw��m�E�p�Z#8�v�`�L�*�����@��C�2�p��BE���ɖ��_�n�J{���J�80��7��G���� T�)`�0$��#��Β�$���.��~��(z�kv��xt��B+�M	�d�H1���s:	���*ڋ�ׯ���8g�0������:��V͚�Qcd}��&���I�E�5 E��s֓0��Э6	�h/��C~����ye(,C��`�KNg0&<3"`��3�.x7X&Yǰu��M�`��G��?�0��mlC ď��km~4���o�?��Y�1fA���<��+�ٽ�M��!�����|?㛴�z� �P0���q����{���f��5�F�D��4F�-C�g���+��C՞�����)k�"�y�[�	f��q�rjj�ƶ3hi�0�d;�/|L��f;��6������P��׳�s�}&�
ת��g[��ߣ#$����}nT3���m�1|�j��8 �o�ӶP �H��]���r��ڑ�d�Ͷ�N��>�����%�e��/H�.7p����P�?bK*��m���D<����C#�l�B�r�0�C�P�PCg�}�������繂�[Rc9z�U�ӡi�����ڡ�4�������vB]�D�p���F���� }�F�Z@F��U���
i 4~�� �U!���H;[��(�L�Q��e�(�_H� s�;JxV����|��~��(ZI!�bgR�jޓ0�<yp> ��Q�Ow?�'O)��v�ܮ�T?�v-�'!��<�>�Q�����~�C��r�jH�%L�N�b�$qm5-�y�$������)��i��)�Yu07�dV�XC�88.���%�	�&��M�W֏��)���&3U�a��o��Z��1x��h���[��5 W�yF]�s&r=���4gk��_�3�?�;�Ä�N�l@?��$�0\�+}/�Y�(aF<�2�B�K���ɗ,�:s�Y"z��ǲ�-�I�F��c�<��"���/��:�c[�i�������z��,�<Th�0juy���j0J��߇m�Ų����~�@���3�[�mm�1��"΅�`]ŋBD�B�D��6�5�n�_��6N���6I����2�L]|�Ł�����t����f��&�t����%���M����0�6��Dq[�K�DLġ�J����K��]"�p����?�}
��,�U���3��0��|G
z6��؇s\Z�yի��Ɛ���˿�h��2�FB�$IC�/ �U��Ue������P\�X^E�ҙ�e�V��t���k��*䟿C��,)�K)���`�k3C��������@���W	�������zW���\3|�J�!�a�uu�f��p�M.�x\�����>����[i'S�#���^�]���\֞3���y��D�3�|�,�
b��=.b��j��~ǵ+`��sa�� oS7Y[��3&i�X�}�h8ںD��ۃ�A�[md�g؆{�-����x,�X���<}���2�$�^�E�i��t��'牧�5���/X����}����~�U��i��@���U^�c�"[���uM���8#O�Գ�"qKn1�.t�
e�7�2�xR�S��q^p��%L�����(-+��%��Ic{���I�e4贯U{#��*�[ϫ��4x���<O��Z�U�P�q�����)�ۮ��!��yyR҂4�&q+P��L�J:�Ә0C����/��������C�!A�E����y��F 3�L���S�У~E|P�J�UDRF��}���:�+;)U�`���M-F���H�;����^���?ܼ7m�����+O�s���Kt���h��aۃ������L��-��y����e	#f���:Hu�>=�LZ��Q���A<���{��<�W�W����L�#\�~���;������b'����q�F��q'���vs���5z��`J �d���+�����L�;��g���U���Zs����%`03�zZW5F�\��I������s��nYvx8s��ʙ�-�S�m*8��Z�*��� �)n�0?9�&i�������]�Nl���������sXcM�:�O����Ns���5�D��*�=�e%҄�0!�\�ֵ�4*|��Qa�X>��ٮ��B$i�½Ƅ
vq��.Z�9�^�ɯ��_�j;�/�_x�Z��>+�m_��Ϡ�]�����ć^=�V�;�t�43�G�r4}�����Y#��'�����yz����;fw��4��-`�JVMÀ�+�U�^��תL�{�^��J:��d�ˀ����ϫ�kvP�HAż?�'�v�4iQ��6֒/p���<����j�Q��v5�u5��uLiz�c�t�3�g�E�����I��:fѥ�
�$MYq�(�z۹n�0���U�+}���'0�Y�4g�s�����3� �K���W�Knq�l��8������x����h���}&`��#����fa��O����*)\0�U9uyb���|���QCO�.���(#O2�%`L�n���Ƣ߲����x�|��w���߇�y�E[g���[��:�A�Q�=N3�;��q�w��ts�e��,ߜ#���0�0��%�
B�.ѿC�x���Lu���=u,���DA#�z��Q�tQm���@B��d�>�RVZ�X����^&�������օW{�5ۡk�l�.����pym����n�#5:{��Y��FN���G��� .<��.�2�R���E��H�k�>�e��Yq���X����� �PH�eG�k]y���_?6T;�-�0p���=��
�UxT�������tϡ���j�8��5h��-�Nm�ڋ[�t�͖C��%�Xb"�_ΘG	�Ǒ����T�U/gp�S��Q���<|5�U�(`L���ӳ�z�k������!���{�V�{˸���D�^� .������ 9���������n}��E��2�/��D/��1�\ey�c�j�$��"\���B'd�嗀�����62�G����
�h��;S�=��L��b?ҁ�!<�� �
z����{|Z�ژ�X�\|��p
���]B�q�R䄟��
�	_z�WV��*`�g)�Qh�(K�l.��z��GL�ڶOA���#}�׶��j�^*��wG��s������C�,+�����+�k�l��V�M�O]*�گ�g��v76����y_��k��sX����#gy}#3I���"f�fz���~{���J��3^f }��o8σ����R��i�ׇ��10�Ҏ�63�~o�M5oy�z�_��7=u�졫o��_�@�7)�`�	/c�lտ��'�FO�U�D����Q�k��&���x~�
���L��p,��D��A�|P問�H6X"Y�$�:��ۥ����K�<�[�i}ע����="��	g�Wnx�}*���S>K����M�����YlMβ��2K$�.>Y�$��4�Z"Q�@H#O�+���Əi � e�����6'�m�h�����-l���g6G�'|ǘ@g�m�I{Y/Zq��m:O=�^=���[���9�G��<��h6}���=d�DN�i�DY�Kl�Z�P#7>�W;�KK4�I�v	�X�����C��Ze�l���l^a����j� bן������hV��C=����_y�{u5������i�o	j��O3�qcD�p_�V����[�ؚ%������3�߸7�V�������d4�1�B�����m���H��� �GC�y������3��8�Ki%�sv�m4/�1���=�
�ZĻ�NyiZ���4/������F�)7����O��P�q�5{��4q�Kj	�e�
:��]$e�y-��/_7���D�`m�j��:�:��ԁ=/���(0J#Qߎ�V�� ���n�9�1^����O67�v ���ی��K%�]!�����?��#̝�?Z�nnN�4��
���w��ʘ�BT��T��hi�ئI��ڶ�B�����R�u�G���cQǏ1h�Hz�5G2�䌚5F���;���E��v�Ц`pY_��������(i5I�~qз���T��4���z��J�(i��*i�|�0���}`����Ѽ���Ͳ�aB�g������;}X�V�����o�������`䩊,�`����B����h�A�`�WBF�o���S 6�|/w��+�V�,�gZ~����[�l�mE����P�,)������a��ۇ���u�[���
�]��������4�3Lȇɿ�AW跫� P�ge��g�̇�E�H��m���k��{�j��R[����[�U|��L��ͽ�,��~i1�A��ne�E�����G�S��'�"��i�a���3{c;�Gh00�#��f�wW�=�"��Z�����lF�i�ka�Ϣ�|���+�~���v\~������shZ.s<���"GK��8�@S�c髞@WZ���q��YzƁK�6C{�-�Fۡ�hkP�y5t0�u�_�V���"�6l���F��=_��9��ĸ��k�|��ea=��������`�ȳ�k_CXy�p��6}���܅��=��f-�zPW#EG��:�O���ċt�ղ���֭�׻��A��~#�d�w�$�ӿm;�E��j�gHܵ?����-d%�v�����~������{��w��%����_U�z��L��K휿��omS�lӽ�;����*����ܜs���ݻwc�ZMFi0dF��Zzy�ޕAK��<���iɸǧ	�����+�t�˰J0	}|.r�U�9H���ǥ%,{�g���r3����y�#~'1%����$£�j;Q��!���i	����)�aO��� b�Tw�bZ��Y4�5��[񊦒�Ԁd���jc�븴�\vH��	�y~���Z�K�v/�zFl�<���1���>��M�H��g��6��7a)X+�W2��@~Wۻ��鏆���]x��x�?���ss���D�1��A<�{���9K�KC#b�BP�-\����?����#���l��Ž�u�ģ�"�^��MM��U��qi�ˣ�r"dF�/`k'�lR���-�G��y�hK^&->Ŧ�)N��� :|�T�qx͊��~_�%aM�;�Yi�W��32i���ϴ�b�����JG?T0o��mB�U��@�唼j7/���~w�//_}\V�ѦAwE���1�^�'��2*�lK�g\�O����[c`G��fnE5�viٿ���`�:�{�v��r��`���+g��o�eZه<���3�V6�7���D1�� )% JB�|�U�R�����i���p���=lS�q�2
�^��4T���
2�)|Z����( VAf�Mx+�������9��M���v�yq.���:�3�/hhD�@�p	$ɸE+�.왛c����b1�LK|]������Z��(\�T���2���1$` �l�߶9ȇJ���o^<k�pX��[�o���"Y��˴c_�(��G����pZ��|O<�[Q/�����q�A��uI�S��ק&../6�؛���3���	3�w_�x�
�6��S�rm�>�V�Ϻ� L����aӺ��v��tQ�dR[����{���XԿ	Q�b�A�HB����vz�p��y�2�\n�Tk�i��1������>a���*�����4�/�Q�.-T�,��V�8�|�<���m�E��w!ԍ��}C�w�f�'��aIa&q�m����7�5q>܆�ӆ�����/#iW�Ͼ`��V~3܆�V|bx2��q|b|Z
���o���~�;v��ϋ;w:Wᵕ��+��!�@pV(���D�#��a�Ad��M/ui~���M}�s��?�?�ް_�>�r���������!��q����֏�J���gBV�~�
����j�T!#����-F۵K΄�4��:���a�-�L����
�a���0������L��>�u����}�8�n���Q�;.�<�V����!KwW�P��2�����2����w�:�jM6�������˫���g0�������cA��sR��w�D"�.� h��6M��<�K$/�WY"y�<dwEyj����}X��^/�]�y��I��0ғ��$0�ey$�Hآz���ͺ�:W�tϥ+�V��hv�}�x���ދ�^����~#-�Cvߎ��Û�)�~|㷑G�Syd��,��yۗ�!�l��O?�}��k�K:�wGy'�H�R��~Nǥ��h?����Ԇ��N^������4\vWn�I�`�J@C�0��?�cG_�nK���B�C�HLC�W�@�t���H��@����`a�в�ʻ��;����d��G~�;�B�|g�{ݷ|�����ϝ�x#��\�uh�Y7p�qw��a�<l��k�.���0�]��y�(����7x!n���(�>�,�$gp_QK$��^�#b�%=?v�uc���a!s����s�SO0��=|��#m=f���	��h?�`��i<l�w}?�|�z��q��tO.ߗ1�"^K���gmSx�$�}�<94l������'��79S��$���~<*d�PA�$v�Zi���	�Y4
Y֣�ڋ��H�Ճ4�ɳv�,��y"J�@�-M�ɰވf>9dՓ���S��h�1�H�9�ش9i���4P�Mҏ���|�_V�)a�`��K�g]�����>:���c{�������6�?a���CSф���96��8��A�M��N3�Ǟ��P>@+��_���}�9�H�����hk��q�����p�V��/^�y�z �'�1�k�Nf��%b��2-��I"1�N����t�WsP]���E�j?�C�o��)�xo1y���?�^�'q
/��`S}Ty
�e�+h'<��n������h �7YO�
r�)�����w2�$J5p���Ǽ�60�M���e��J��6�ݳM����֪]~��  �IDATǻڵ�>a,���Z��Z�mZ6?�b�Xoa��Bv�|�n���$'~Zx
[#�y�:����g���2�?����I7.p����r���˳l�=�ki��8���f��	_�e�hu�I���g3�L��AoVpۿL|���珈[|��c�i-`R� +@��v�W�曢��_����˜;,�D�����;��I�uze[��-���1Gĳ�AM,	�ڦ� �ŏx2�� ��W<sC�ψO����p�.���խ��1�Ov�ɧ(OZ�Ü���B��Zi�/��=�����6���!L]�B����hi����pXc�SXi��m�s��~����a�<���S���E���H�����f���g�f��i8-���fw�I��O��(O�s,|�Xe�^q�-�g�-�7R�\��G^�NݻuW��~{��A����G�?���ۦ^��?�cM��z7^�O���6�xEZ	�D~ɋOɗ�&��~+-h<MM�<�c�vܷ�?}|��)���0K��֍9��lê���~5uba8��,#�5�cj,���M���<��΀�������9$�����Ƨ̞�^"t��|0�\���8� �t>�2x�y��߄c.���E���L��ߧo|�`>���ٹZ�a��;�HϣtX���E��D<̎�N߱��d�qp�u�8��k�c����6@� ����Cf�01�=Z �m�u'�kĺ�z��{�����ydgM�[<F�r�M7<��N-ރ���l��l��Me�l���lWh�V�v�sx����X��ۀ����giav:� ����́]��6�<�w����'͙�KH���Iέ���ZO>$/�?f��%����E��	`�m��Eڷ�<��hӇ�����_���ү�	ڥ�M���\U7�[�t��3ݶ�Α^��	�F�!P�f�p�)�<8�H]/P�0��<V�g�Y}����Z��֯Y:v�x���/��w�)�"L���^i�]�L�cvi� �Bڱ� ��78ut��,[L/���,�����pX��&q�>5}�y�aw���G�1�9m[�L�yƠpɟZ^$|��4^}]z��C{��<.ۓ4�㻎I��|���I��<ϭp l�?�i{O���cЃνky��?T�k?;��C�*�N���z���W�3FX����B �E�}��������F"v�>iLh'�*�+�a\��1�2�?�ۿG�e�w�I���H+�ٶ�i��k�.��7_��q�'�&�ه�"4��s�8��+��͛����Q�겈'T����-}ˬs���b�i5�Ai2�-;��D�A�8m ���̺�2[ּw ���a���	Ÿ��op'gW�+]����� �?W�w��
Cإ����U�����4ӫ��$DN�\��q�BG??�=(�ph�����ap^'@x����[��������}�:vmS���f��@�d���Akz��߯+���Knfi�9�I�tJ��*�ku�8)����Y� \����xt�n������k `@#�� ��y[�y��<�e��h��Q�τ�������<�&_�v���<�+ÝZ �,�o���5��q���|�Q.D��!d\vB��~4�?� !8p�eCH�iL�5�{;�Cbh1E�&�}Y�'p���E���143����~F�;�ot���|���z�rj�b�Y=y��#+��`�j���IN[�xsZxډ���w�o�*ڕ6�*MZK�K���E����¸�tq��$�q|�-�g0����(�5"[�Ĳ�i�[j.��؆��p��1��%��c�slWF�uO��~���W�3���M�N�`�g�)l��#�������9��#��N<c���7�h��[~��٦5�f�pcg��Kg�&C�w��J~�p�lSC]�+Ǳ�7����X�uݱ&�\i���E���p�����ކO�4�Ar��~P�H�<�!E�t�/����=��1f�X�kW�m[[$�ˈ4�<��<��U4��5q��묓��n����ƛ�$��j�,��e��k[��(w�k{{��K���)�.�u�a��|"#��d%H|���0	0�5{���M1k�Ⴐ%��-GDx(գ�OО,�UY��3��-7K��$R�O������'j�Ŝe1��Z)3	�c�"����(�tb1��Ӳ����T`ې�4QO��<��I��$N� �r,�s:���]��3朹��x�z�f�"����4Gw9;�m�iV=@ϘGLӡ�<��yu_�]�bm�����R�k|f�vFj���E������9Hw�e>W#�+�U���H�j����h6&��LP�	^�6��L��}����䃗͉G�����ٖ��f4���0�A@�r�H�[�$�W-�l�=ݬ]>߬_<�l�P�4���&���)�S;Cx�(����A�h�f��W�f^7k3�������2�c�<N��W̠���;U�l8��{�9�DB�[h��H=̀�G���֙�f��l��0ۼ>ò��٢~۩)&�Z�>�88p���nCg����j�'�����M"HmN1˛!�I��o���������f��h6��Q1C����XN�����c��@�f]z���<M=��ӳ,}�۩ڕ�3����	Yc�3'e�#����ta_kiC�?�00Fe����G��G{S"��<�>eMs�'b������W96�%%��F�����cZ�u�~�w����'?j���72��!DS���Ǒ+����F��~cm[����;�
��/�X���{�<N�įp��y��b�>���4�L������q'�3i8�#�h��4�+˱2!v�&'�b��dG۵p��b]��G�~�qs�Ӯ>hS�>I�w�u�1�(���C�Xl�]    IEND�B`�PK   ��V*�.�  �     jsons/user_defined.json��]O�0F�J��Ċ��w���@��v3US�8`)���UU��Ja
�vi�y��g�]�����?K]�K�_ڷ��p������r��`�c\\�q6�t��b�ʾ�!��N�8�I�-`�#vS��LU&x��SD��(4�YUfU�aͤ
���qt��^?��u��i�C��r_������	s���r`����m�b�ru�%����z>����#�!#T���$�5w}h`/�u�M����5c�KS�� �8%(�DQ�=����0{�g]H=��`��F�Wh��*������$���3��W96�s}0����C��Ѿ3.�N(gg����okU.VS�CHd�<VR��JƂk��c��������0�B�韀G���AA�`��	��@���9
��)�K�����l"�=��i<���'�'�1l��PK   ��VZ���=%  ;�            ��    cirkitFile.jsonPK   ��V5���� � /           ��j%  images/1198b7a7-cbce-4bfb-9393-e70c622bc3b2.pngPK   ��V�<�ѵ n� /           ��w images/b6c897d6-7294-4140-aae4-5fd8f682e5bc.pngPK   ��V*�.�  �             ���� jsons/user_defined.jsonPK      <  ��   